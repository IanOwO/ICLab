`ifdef RTL
    `define CYCLE_TIME 3.4
	`define RTL_GATE
`elsif GATE
    `define CYCLE_TIME 3.4
	`define RTL_GATE
`elsif CHIP
    `define CYCLE_TIME 3.4
    `define CHIP_POST 
`elsif POST
    `define CYCLE_TIME 3.4
    `define CHIP_POST 
`endif

    `define CYCLE_TIME 3.4

`ifdef FUNC
`define PAT_NUM 828
`define MAX_WAIT_READY_CYCLE 2000
`endif
`ifdef PERF
`define PAT_NUM 828
`define MAX_WAIT_READY_CYCLE 100000
`endif


`include "../00_TESTBED/MEM_MAP_define.v"
`include "../00_TESTBED/pseudo_DRAM_data.v"
`include "../00_TESTBED/pseudo_DRAM_inst.v"

module PATTERN(
    			clk,
			  rst_n,
		   IO_stall,


         awid_s_inf,
       awaddr_s_inf,
       awsize_s_inf,
      awburst_s_inf,
        awlen_s_inf,
      awvalid_s_inf,
      awready_s_inf,
                    
        wdata_s_inf,
        wlast_s_inf,
       wvalid_s_inf,
       wready_s_inf,
                    
          bid_s_inf,
        bresp_s_inf,
       bvalid_s_inf,
       bready_s_inf,
                    
         arid_s_inf,
       araddr_s_inf,
        arlen_s_inf,
       arsize_s_inf,
      arburst_s_inf,
      arvalid_s_inf,
                    
      arready_s_inf, 
          rid_s_inf,
        rdata_s_inf,
        rresp_s_inf,
        rlast_s_inf,
       rvalid_s_inf,
       rready_s_inf 
    );


`protected
;ZEEF6899U/(WY+G1QR.#SYW:IaH[HWZHSd2(8<dbR>TMQ8Fe.[E&)/D)GW/AMB_
A-AW1UBg]P#0[dJgWA(QH2=F/Z+SaUMfGHf[1V_d-=GLaA6&UD\8:_JNH7?9/BBA
/E6[QZWA3,7Bd;I[^/ZAg(>&9Kc>)C9S19+/PD#Q^(aB9QX8-eSVI0,1cf+_5T&K
0HdA.HT+C..eHd378F7WB2&S?(S5b2;TG&6II-WfKNb^C-B->=\PW?dZ7F.>5H3O
5ES,[,0egZKDb)H&ZW9T(^3Lb?=U(VONcV9fEUF/;IVKKOB4f,gDE71\4?YTQ88D
TB,M,e;f?L^?A#:BMH8+#/1M8,e4P+/O;L;YG0OH@K#3#+&K8.;;O?Z:FDg7DTL4
UM(ONYCB-Ve;E5?La+(&@/KCK&W+\WZ=;$
`endprotected
output reg			  clk,rst_n;
input				IO_stall;


`protected
_b?X&bDQFJ;B2W=VESfC6dNe<]N;86NA_R-/IXQI1Pe/[>e\IC,</)&9[fU8dAO^
D/>>X\3IGag0Q9fM<RTX1XP?#J[QG2^LD/ABJ+.I5Xb/F$
`endprotected
input wire [WRIT_NUMBER * ID_WIDTH-1:0]        awid_s_inf;
input wire [WRIT_NUMBER * ADDR_WIDTH-1:0]    awaddr_s_inf;
input wire [WRIT_NUMBER * 3 -1:0]            awsize_s_inf;
input wire [WRIT_NUMBER * 2 -1:0]           awburst_s_inf;
input wire [WRIT_NUMBER * 7 -1:0]             awlen_s_inf;
input wire [WRIT_NUMBER-1:0]                awvalid_s_inf;
output wire [WRIT_NUMBER-1:0]               awready_s_inf;

`protected
SVUEQeaXTO.-L/,VeORQ]+&?]b#RN#0S-1/?#@Gg,7PgPZ85a,ae()LBJD4,7-7-
fE]@=&\(6=dG[6C-AeU55COL4]R&WZRP(5W_O#\]L=TgC$
`endprotected
input wire [WRIT_NUMBER * DATA_WIDTH-1:0]     wdata_s_inf;
input wire [WRIT_NUMBER-1:0]                  wlast_s_inf;
input wire [WRIT_NUMBER-1:0]                 wvalid_s_inf;
output wire [WRIT_NUMBER-1:0]                wready_s_inf;

`protected
d;Cg?2723(Z3=/KS6-XH)GBe:J,BT_ZfA961Z<;@VB;4[)F;ZY@75)Q5L:Vf1[5?
\[Qg4g:@-/b-fMf4#G?A,\G+gFST);IROb5+3DTWb.,4F$
`endprotected
output wire [WRIT_NUMBER * ID_WIDTH-1:0]         bid_s_inf;
output wire [WRIT_NUMBER * 2 -1:0]             bresp_s_inf;
output wire [WRIT_NUMBER-1:0]             	  bvalid_s_inf;
input wire [WRIT_NUMBER-1:0]                  bready_s_inf;

`protected
8N[C]82Z/>\Be82UgOKB:0c52R>W(<g@FI9.JF,:G]UPaa35E.6T-);KYKb/(f&)
_/#5TgDHe@_CJ>(c^#;AWa.[.]+X+Pb2Q>S,eM5>5fRLe><efF?XC-C/bZ@3^-DK
@\A)FTHYR5H)6PZCD12MW_.[6$
`endprotected
input wire [DRAM_NUMBER * ID_WIDTH-1:0]       arid_s_inf;
input wire [DRAM_NUMBER * ADDR_WIDTH-1:0]   araddr_s_inf;
input wire [DRAM_NUMBER * 7 -1:0]            arlen_s_inf;
input wire [DRAM_NUMBER * 3 -1:0]           arsize_s_inf;
input wire [DRAM_NUMBER * 2 -1:0]          arburst_s_inf;
input wire [DRAM_NUMBER-1:0]               arvalid_s_inf;
output wire [DRAM_NUMBER-1:0]              arready_s_inf;

`protected
^/I>,NYPX8XNH>eQ3PYCIO)?C3EA@M;UG0]MS6ZNP7[/aEN(1V6R2)BR_1&BOLQC
\+ST;fM9Xe&#B-AHIbB#L4Z01_R&2A\@JNTR,@UEf-C^@=M^:H85ebK<KAYM_c;;
JR3f89fC;+/,&+aI\cFe\BZ03$
`endprotected
output wire [DRAM_NUMBER * ID_WIDTH-1:0]         rid_s_inf;
output wire [DRAM_NUMBER * DATA_WIDTH-1:0]     rdata_s_inf;
output wire [DRAM_NUMBER * 2 -1:0]             rresp_s_inf;
output wire [DRAM_NUMBER-1:0]                  rlast_s_inf;
output wire [DRAM_NUMBER-1:0]                 rvalid_s_inf;
input wire [DRAM_NUMBER-1:0]                  rready_s_inf;

`protected
3X[gOJ9QI7fg^MVX^4dU:EJHHTENQAe(b&.&SERRe#1L1ELR&/QV6)G+)QSg8=0H
-[]?:&>gLeaS\I#1Jcc)4\TeB_QV1[2=_^-R+4]-=4_<<U@Ge/(aG,:P<</VH/I\
bA,Ib/.+-#dc@f1bY=0S&/5#Z(E6e;5,J4^O.1bEB<HPb?7/T&>g\g:58_Y1&<f(
g>Cb3HQ??ZPY#0=6:\RMAc/A[Tc1E32W5?^H03]//\S6&5=6&-1(gg1bK5E+#LEF
)\VK];aUdb2/e\&.>U<+OTgL8(7g_,=NZQ[U,1NRaP;3QfTVg^=SI)7)L^VcGB;T
U>;.HQ,8cCf;XC_SCXK,W,)c?-YdK.5>^\>CEF[HLXC>1&4bc3<J@&Ag,M5YM^/a
EX0f:Z6-cULS[GdO^ML:+H>25FI\MYI[?@f4S/0)&>NL35<,MNRFO4TbLdLU.:PK
/6fXEPFZ<W9VZ,;a71OVX0SU&3TP),LZ<VI5#=)SO0I28Z-VL;A>U@6\Sd2]0gU3
PAB)GYgRY=b(dT?718&abL4WG@_S[]P0=5>)aQUGE8aQZQ6O(+1KRP2SV\8#Q[HU
\#=2R&8b@9-e52TgMG-WWf\2g&S6)&6WKME9(U0Y64<f<EggXAGYXO@1SB1/[JdV
c5BK+V8Ub4BL#E[c0&PTO422KB-4e+IO&U(JK_aZd-g1V+;1=?9LDHU4##(B-Z8\
DHPD0F>Y<?EKNPVL^_GU,VK;W<dN7IQPU_fZKGS[8(K5L=.bOb(5V8B#JKC5_&:D
97OL^d8Md^N-I:J<6+6H7fIcF)8<Q1IU+3_O8RJY[#5YOT>G1Ve7f&=INULcRUZ\
R\KMEfT.PcV@TAC;+f63I/;RE,EW72Y_]gaP]39/0O.H15I]/=;AV]R#Z]]fGH0E
;HbYSOXQ:/<BD.CP39>(NNe]gR<?=7GZ^OEZ)V6@]Z?#_)U>-LgN=85PUO4Y6_JR
65/f#&R(]NT=JOHA]b.agPcD;F8<2bW@\]U=]Pa5:L)PY-IZ(:4Qg[K-R05,N-<_
FLOF7a995,_Lc>a=ZdV84N50V[RP^_fMIB8#>d3c?bQ<Q[J+(JNMb&3a@b=-[P#B
JNGN(V2UB/gC+X,WdU<3500EC<6cN:Oe#Xe9WZ7LA(EE0M1@1CHf]R_,4cD0d0CE
++@HZ-M:99(T-f&7B\>@\[C.N6R;>3;8PZfaR5gg(c\XYJNaFd,(,6>//;RP0IA4
9Y1K+&=<XK0A]LAS4X\f-a;XT@9VL9ObP>b\-L]a)XSPcZ)4@]?AfDU6Z=);d.KG
RM(-,,KAFG+P24a5A.7b@cMN?T2(NU342d?;g20[>38VA>c=0>XLA&[&NTWCNVD.
4+U:Mc>MN5FW^8JBe[KCe<[O&UFPRAVH^eAS_IR]Z^P/Q\1.gaD4EC84S4=KH>Z\
5ac^G3@50([QKc^[715<(],4=^T_>#FS=[^F9PQQaLH@O[;J[)a\V7Y7J>RD>H[U
9^UI/)YEKGIV2[F1FI5)5f-7(g0C^Ga:_Dc#eHd^QgA9G<[<JU^BFY2T.R1Va;@4
2=B?2c[T9E1KGFXg6/K,;^1.5c(&cERZe^7b;Sd4JFD2[#-gTVeY/WB>G/gF:UMP
c-)DDZ)BZ,@;K/ZWJ2@EWD&6Z>CeO9H@Z6<QFRd/GP^:J\D<UGcDO39Cdg)-(eRU
]MJ8,R8YIG]_81CLBaPSH-[SNa4_L]V9ESC/VB#UN^1bCT7:<eP:)::M-_3M4)\^
IVQ][P1VBGf)7-/&HX?&bSUABR((e_H>C8ceGR,N+GWG88YH:E\&65W]_&6aX8UC
9W<\fBK8ZX;Z;(PY[=_NAT+#/;_TaDP97/T/1]#+GET?_Ja;/A(d][<GF90<d--8
CMNgH5aQbXJ=^C.Ma=(V00@#4MI+b332S<.BJ>UL7f=YKfaTZZb(?<\8W3ES+fgg
<[D?TJ28:CJ=WBZZTG76c8I0>5R459Df3>Gcf,UM;^2:_Z)8+.@@+LHT,X^.,G)<
(17\131EceV^^>K]gG/E^GL2?J-V[W64cW>#(+7LDLX.FY,Rg&_\Z<L\9e1+YAA;
DWEE)>QNM=ZLdR?OYR:MNCHW0^&B7dAa4O53[D-Be@9+TJ+GAc3fD]9#J-W.WEa;
HDPXVLS@_YZba,D)c+_X#5d[cF5aI=D_82-K?]S/AUD0M7;NT;F#;U,-+ITcR7Gg
g(F9V+\7DZ9S:;ZO,4W[,KO&284>6&_VX&gR/N&S2OGF\:FaGMKSQ8&VSa.U]-Gg
+Q<KI.6a[f/0LOd;D8L7QH0OQI_]_BX8Q;DP##UQaYc(<bY#@])_@0=J0FBA,He=
.R81B^g&_OSMI5HY14^T@[-C63GBe.^@E?7O\H61ICLCe[&=NDTK9HAP\gQL([3J
G65-QJO(0b\Y99?T388U?AI,I],>6a?Df\/P33KHR9=19Z6SGcJ>1dFO6PYA@#U^
d:2WK&(USU3?-2M3MfUBf,AOS3HLA<\MRb@TSQ99MfSb^1M[Y:[)e4-G]O/LeB]6
DAR2FEQc<M),AaL_]A?>cBX^ET9L-TWX2:^9;S)JY0aC^bTKV:Zb7JAI5eEdbO5D
+[BQg(2I,g/VV>?Ag;)?Me,?A,KL8HUeNf519_F;&,;G1,gH7:>57Mc&Lb+:[^Xc
EP-^^O,YY<Kg&T]SS&@XUR8T\fcD?K5f+MFf)1DBXT@YA.Sd[.A0aU.CD]72MT.(
(\)8cW-B-W,5GgU:FKM9T1F7L<e/4@c8A&?G3172T4RCfPH&RaI#FJJ5+b@1=TIO
O=A)E6Y+4Eg(+\_Y#\B40EB0HgLa9d1=FLZE?AJKdeCgN)IDX/FXB3LbY/dEI#V&
[(?CQbbdP#GXfW/B;414HXe93IWLa;-1UQH-PC<:[a7U=]C-IR,9C&&[ZV?N_]SP
;2)<_DdAQZ_-SPDZH:D37G,+XOFW=Q#KOA[,6_GO>U9ZAS,RV3I#)J-(KELEUJ2#
I\U64#ZJ6BRKXEOUf_&NJ00X@]TB\WCWCgd33@9E<XbVXAIG0c4Ee)7;=R0(R.^)
#R#M8L.5?AKKP:@&#=ZB;=EG16/8=V;J1Q5:44OeF4bT8;XV)TaQ8+O2AHg82dSK
U^SF,#3\IJgBN81KLHDD.XOc0U];Y;Q9c2L]EaQ#;GJ&Y:KSWVOJ^2.OPG/KI9)E
P_XX]=DGg8CG1G3S,+_aW.#]U93bAK7N76^ed-E&I]Q=,V9<XW^>:&LP_O_C:699
1&O2T2@B\H9?;OAZ/J6:&_YJTT(M[?2_J0=U:[1M52+6ef:dI_#/79;W3=/Q[0aS
@0OK^R5Gf):WW/ANDPZeOL<F9ZLTAHRLa)B6ge=;(.8+W,CQg9?@11B)W9KIE5g6
7A.^95#Q-f0X5#4N+?2\0[).]DA_2Y)8/>4:bgM0QM>6f-./_f&W.dV;/-A1dG\B
1<[)36CQ.A_@>1\FaSQ]1Q\>5FW]S=(D:#@(\N<YV\:]f(@]Eae9,7fJe.-d3Y0e
>N=:fY_@G2YEaIF:c4/#@JaBRJUA4]9?L<Ra\8b:fNB4#dZ\9(?8(\<\VY2\^>25
J7a-^5;Y,G7e;EOaF^9^161S>0D_#B.^J6BO-H=8Q1I5^:W),W81/YEI#;a6U+?X
GV33:/Wc#NWaLUG/I2aM+(_9?&(1[J+2^L,UYNJCX&NL2+De-BN+QaRIb+,:#;]C
_EV\gK&ZH.WeV]QdOIM#ETIb&UB0CDT5fMQW7e38<O^RIEReD[6+HfE+,]ca0@Nf
8:/5ET1S&5C\?IfP3L>@2L]-;^LR&HE>SaYeH@D+.O3]/+_7X[?=\^#1..S9]\[7
]3E(HfHf&55(CX0B<fA5O\b;eV>?\E.]-O3(SQ.SEE1Z9:cbfeP3=+DOWF(#4\H5
d<S9<\2?3-F/]^ONeeW3SL_C0_APSafLQ=DUCO9Xa>F4E-L0eB)1H#:\#3@C\\SP
+U<VFNW:#Na_X<V;M7+KbF)gRG[4+5fKH3[.OgBZY.1TD\e+)(T=HI7b2EU19;4.
KIL;,JS/\<]P+J\MOYRbZe&.MaZ:)G62S)ZNRCc&gO>XLQ[F8dVJ=E4:0X3<>)B-
:L88N-;S\eDGBHYT4N+,/6#&R\Y/ENZ\_GIEgIJF@[M_2\Qc=OWPf4cQC_NVCQQQ
IKR5CJ+c1TVP1J7JM^#_Je^S<)1YfZ8LLdaUgLT,dbe=?K&&<gBgBa>Y;NK6FD.0
]J;I0L?HfKH2I^(4PX])=^bX(Oa2=O:=[3RL.[N+0RP:JO\D_dR9VC+&13_2e2_D
de8QI)VdX<#\VA@aY2LUJbYO)H+f@-:+WTE,IaH,6C&8WAZPOXC_CKaF]JOaL]OU
fQ.P,OLVaP?;I\YaEfA64X+#8[OKFf_+#,I=eV)T\:9]_O#Cd6/ae+&fM\LM;=#J
6<<@AW-:S3F]KMNWQNE0&:c:IdQbUT,PVZ-VG8=[3F:.a36-eQ+/D84IGA961]C3
G4c0D2\,F?X#73_C(.UP_]Tb>:T>(,;AEaXLDFPG]XRGCF<\51;ZS(F[3GEc6DHK
=?D9P@<\W-DQ#(-J&>283_Cdb:=VFZS&QPEf8B1126L@UJUI=HF^B)?,-e9>T<7.
E59G80^_\a5-?[=,]G#aB+ON>;PZO3)US^23A3?=FJ,76X[3eUSY4(F6VJ:eRRdC
A?9L?29JX/A3O2&+]c=FU.Y6GM1>O5(6KUYVI@W.Xbg8dD^F8)]U3gKMZT+b[LL:
NTaX2U^^c:K,L#&,CEAg:SfWW,_@<d8+)2Z^S]_?+T?[[YAHHIU6.:f19\?O9M&S
R(@AG+,@Q.>CJ<I^@=T^OV1>9V,.U1(/WS<-Q05VO[K38:4^R718V0\#26^RQDW_
JU97faR<AUP_QN4]G7fIgg7J142[]^7C6C4N^:X9Of4A#UFB\eRQ/CGgb#,O=EM/
@I)0J[+6LNQ\0_(MDXRW?5S>Q;.GHOTUU6LdD@Z:_1P(FV/DPBV2]MCD0F^O[3Rf
Zb1.0TO[S[d9L83Eb[)0fg:d6[IHZTNVX:5H+^\V#D=K330e-TEe?L.\RVVb[YGZ
FD[74VHHM7VM,(/^U5JbCe^7f[54(d6ZO@(a5(XdNX4+D(#,a6FGO5PP46J@?AV/
_@,Q.\EB6YFf1GL4Q-X>bC=1?=7R]\4eFJPN-HF]^_A<C@.0+T9-5=[cMEM/G,KV
)dUb5]fYbXK@)g^[;cG9=b3S5b1QLZV6#WQP@7@;MS^-/TYbG5NR5<b7]&W&6]QB
<S:[\-780,TbDJOgaM5DgeZI[Yf2E(3S](Zcg8M[W(;DaO[9]93gE?2d[;-P0+_3
[F\L2&(ANYa6c&bB:-M)\d>Qe?\,TL&]TKHRQdU<FQ77b=J6112R.);Xaa-/@:cU
?;=2#7DQ2HV&0TO]c6Q_R5W;U3?8D/85/Z4.=W6bC\O\e@,5)R>&@L9A-S0AEEJd
@-]fdKA=J>#>3^+AB@:Kd8C_U0-C^CZD0]6?JJ;d13KR#LBE23#Q.RfGI7Jf[@:4
Y,J2GEa[ZYAEM?D)a54edQT>O)N9A,>]:W0LLIO.T,#,4b77[Uf/7UgS8(1cFVTC
:Z4f@-MPG<CHI6@36Z+&4[&-2E&e@21_7J=DdL[>GQPc_NT@,>B0)Y\XW6&c5S2g
QA2PBfV2:JP_YSa(P,LU0CK=-RI]FJY&g+)V=R7Y;26/H[9Y]C\AW23eAAJ>X-Fc
5=V<ZFH>,W98L(JM/K@/_@;WSd)5)QRd[6@CMRA;T>5J):e_=;&N?2#PW4++C,0P
=MUG<=.&9UMfRLgf0P:DW>STJ^VEd:dC[TW7eac^<Xa0?X8Z8U8a[:g^6]/==YB1
MB)Q[ZYgcV&_BQ1^[GS3K,]P-66]JM&Fb<US+a03I.QIC+\WUY(^5Cd=-:J1VQ)Z
WgA?-LZSLA)Z.Q[3UL[a2gH05W/6d)b06D(HJU\a]g:P8:>),50)fSIA9V\.(eN4
P:.KAIeEg.eY[F/[=.da,I_#@DZUQBcESbZ1[F..C_@c?H<&K\X7D[XP+P/(3KRW
.@Eb;]V)-fR-N^d.Hbc2g#b[T@,.DJZ6RXV594476;.aAfd<<2J>HB]^->@G]^d)
^F9U)^UPD357_c(QVTR#U-3;LF/\,Ug#^0KMeM1J#5\D:I;JFT98X1QX)LA8[5>I
9_D6)5Fe+&J_LZ4S_[aN9N?:?L[@,,](b=7Kbf]Bb3=G/643KMG9WdH=8K.HCU^_
g(6J1P<&@056>RP1c-YgGXOd8,IT-JJB8O;Ka]+6,f(7JNQ6Y?Dg6<eVDWO1Z)<O
QXf-MS^AfXGP=?7>?Y0@@D,;R_1LWLDDb,9B,60OQa[5?Cg>:HRBIV-^d<(,WE2O
8C-MT.4fQP.B/^DdW=gcO>/)1b77[#;)7K0ae@f>3QB51N/0Q/9BG&_-PNGf<4,c
]M[4C]a@3aS7EC-2Y84fR^Pb,)Gf&H@[_:A)M_3Ig@(^aPXS)?R\[/9HUF^&bZ=N
8^R-D08VN2\UUKReFWJVJa5:AE)+3K6;ccT>;]K,ZF/c1e@8_(a/]TF0BVLM@0YL
4PTES2?g+96b2+P5XIB:1Z&46[X/G[3OcY,8W-NG+8a>0WQV)eTQ=(F\Oa06;9g(
&THOcGM;9d:FeI2b;gJW[+GG_b9T/MccEB]5[Tb>G+,L-4,0c2I/Q]0<Q8A.(OfE
cHe-g1N5dUFK9H65Ue2G?ZENd:R2:^3GY+:5=#7bVY_1_e)\GH<J.,>JMDV=(0D4
1&9Tb0UCAW^Z<S2_+^^QdL6,&A2JL,S+?Sd(#](EVZZN&Ag/3IT+CZBYb.1<Kg,#
g?&UJ::R?>E6S(@0O-Y,3UdP7gD5ON^[-T\^(B)\)JN=Be4Sc4Z=BX;O^XWE[:A,
G29K85J(De-C&LDSSP([Ke8_@bD;2eCV2DX^00AP.W^NRU/,a_U?^K4DSf6W>><V
0MO^_A)Y+,9AV/HB6#B=G@6EbF7F9LB1Sd+W&9Bg[/)7Y\)R)<H4?))Gc9A]0>d0
M44V/+X>TH:7BUX738BgLS1K?O.Z5OgCG(=PXVXH_7?>@Y+QZ,7B/7g7d4.Ze?dc
fAPD1HTV5IB@Of.86=5Z:.d-8NcSe>e@-b1#XCJ&:9<#(#([2^HE_Q(FWg1)(/G=
,(2RBRG=FM\LA^19Zc7[V5QO9WZQHBCY@f:6cR5:V+38YeRE=@\KF5aW/NSc[Kd2
^cf,P&+E7IgF.8f@Zb.6[.ZB2gI@.UBcL4b5OY)T5JVEJfQNJ3(1(JP=9eS+Q+AC
fF8/,FIMB7=Dg.AGfcQ#C9.BU8[,eJQ\SRbZ7_EU9MX)W4I2PaNU2^<f+#A94^6+
e_06=Je(.)JW/NP^7dP5-&#2\?LW&dfeNAU@=3f?#CNOgJ;RUU5KF2Q6T0_W,EIR
OB4Z7ZR]D==XTPf.aaeK/?#A;:R1B;>7AU11=Z1=:23E96BTM3J5_A-_]]EMg59G
)HJ9#@O0H;=+R&#UJ5V1g7gNdacNF).OeZE=L]PM)=H6D6Y1d/\.JB\dPNIWDX1,
Q<(EM/Ug+7;OK-QJOb#/;QA5@M)eITgK_T_BIFGe-NUC,KDG;g1&#K?1C2Z4HY;^
J_gd):a8=0bKYNdT&d@]2fcNR.VRY?TR>\faA>@R2E^Pe2A67;C6,KWKM[9=S(N@
5)#/[RYYHDF<@:0=F,KKT8GE-;//5/IBY6LM,cNF?FP9Z=E0L^P36f9+fEB+P\CU
A8dD.D+K./KdL@e.NJ@cNR^1[_FgED9aPf2>Hg4KE:-cNG9&g0acW04;TZK)1a<:
,<+<YG;V>)G-b].V2VI\7\3M625JOEZTDFI:NKK3GD>Ead&^E>B.Yd.^7CX\-_a4
,R=+3CJ?VWXC#>-#\:Dg@82U,_Pc0)3YPEf12H<.-#7?RIUU7/8WXf2MfU.V2O;-
KN2/&M@/5Z\+S0Ke<fH<&VE.+66BRHeW<;)I^b&a_9@\1L69(_C:<?+0:WSQ#OF-
2Q.:0HV2\T8<&UC;@L=BfS;8EGJ>KB;)fXI^RR+gF2M9Hg?D:7N7S3[7+=H0)U(O
]g5^&UZ+P9ARQCb#4.[4-[5^MZNdfLRPCZI2JIHcB>3F?YV1.4HT5W7ON@PdPHX&
+;\Z:<beH/Q&/FJP)2UJ0&L9/_d[BPTJcf8IB:IFb#=4c29C)@JE_CAe:b(#7(GT
#YZJ]\Q1_0=6fbQ)0(8#>11aWD/^c#PaF4)#AY>8PZPE#>2UX-4/=28NYd)WQXI)
X<N=^C3UO1B2O77ePKbOL2a@KVf4V#=^C:C[U=(+-c2[D/])W>OcNQ5[V++[Q07J
c</9QXa.5O&,Vb8_:bSMd3LQ>J3N5,&bMD1U28[L)AL724@7).RO8<]0DdQMY:6T
MOceOV;E^L?7_Z.>#b<@:/<YN#c__VGJ2N=d,,=R:c4B5?6R&(Lg?-ZW2W;U6#44
:YP18+7T341ME8Q-,c&>^JEDX[T8cKe.N\UA[b8UbaALDEPcB(bQC[C1A6EMED?1
SgCNS-@&f_g\.]EKge]&?;-ZeT/B6QFG&-JBL.Bgf&(+;/7g.Qb7;3BfR;_Q8@5M
#D;K8=WVEMP(,2_79<,S^&_B4#<2)EI;0e+[4dYHTdbQcE[gQ=LD:B\OT:8J4:O3
UCC?2K(aQE1LYW^^]V;=I0WRMXcIE#F(JXSa(g6QWFSR0g8bgJK<Fa;9^&8bM=NH
:,J5&AKPb2D5>@9;edFM>VYU-NOdDEPKZ6792e\.6B=@cNW1H,118@WA[<=59,4A
;KCCQc,84C[HFeP2cNePXC5(g#8.(H:+cK[#M)_gR.K:NMV]U/gPV4#a@#E3Z_3-
^Y9Nd3Q6BSIbTe^Qg/#8P;GK:K>,APca]D@H>#/4.49bTV45<O<b&P^fGB01ZLaO
:BMN5/#_^#\[4b7eeAHT0Pad?gTdR(ZJaR+=,;.#aIc9aO&AK,c_Z&.M&Y:.M+R>
AK]Hbc>3?+@b6cb=26dLg7Q.UHVQ;R.DN(0gFKBKY[9J_fNA2?:9R/=K(_>CVPAO
L@OfMX7L#ALa;VXCb(W3?NKOUDcfd4RMDAXKTN,[RCN#7[QYaKAQCSPEa]29:+8P
K_,.<@2UZY@1FEM+J-13dMV.1H7gALVS26Aa95b9VFQB.dN?c1VZ<Z>U#aG^:HB&
)\S<Q7[XKV4#.@Z.a;@P]V0(7/PbcU<RH5bU/JN\CC-/>IA9PL-\WW^P>ACD,ReP
cM+WU-a2Ye6LUDBS#([T1cX7PYTB8BR)Q]gcJ3f+McR=QB=O+=[VQeSg-9e[<#+-
4/g(A^GHXBC\0-7XA];]QA34DBO#/P@eTgI5I,6dH1SUJLE&PPLE52?MbO&a(Y:X
ScWfd]Rc>:4<VABAEF1#/NVbBbeS[MPYF/3V9(_c(aIM:R9WGc8]3X=W,D/4/C3d
3B5+;]#6J3?3J@ec=CBJWFZQ_:VZT540d-0N8,+2?aZ^FA)?]-^PQP64BN8g\f\g
FG<<-RX<[D5).^BL5BVSRDgb)\0KC3.9Q2FRQJL8QC[>d;PA#X4\(\DWeM=,P1&C
LW3Z5N]UHcN++_#U3&V]e82C>U&,)3U3Q0JV8A)^/94NMdS(Qf33U5&ERUILACf2
^f]B6bHaG#3>.DN7GL66OF19_Ofe2EE^bYgQ#X)3^[[QcT8S2eb<+#IINLGA:dUI
ZWAc.Z&dLIRX7IN,T<-TG@W9\W=T4S<KN:b05Kb89g^4.3PQS#NaIROY/PFZ^2Aa
Wa-I77^\B49;U;N5_CgN&>ANcPLA-UY/9:]J2CX0/A(Z35)?]97&^#72^QMQ0()S
XPF<^UJPFA5<V4Rf3gIIg2_0K-L^7D2WSU]8U8E/.^PJ>BLa;0O&a<=ScLPBLJ[#
.Gc3>OYHL<K0YKX&&EGNX=GM;(ZFeGPc@9>Z:]I3SLT727+GW-#EU#2<Zec?]c5]
\FQJNDfCOQ.#2)>)0\c_M=RLG-KYb99,cd?Z]/[gXdMK\.7f4[H12CY5K(;a7B:A
ESBG30Bg@]/fZ[^CE4O[e9=^GcP6M3gG3-dWV&K+JLOY0J5[XdeUF9N4dJ<BRK#)
W53aeY-b@WaX+2BOZMa7^O@Wd05E(^g_;#-EGY^+\60&J;:GCTV#4<D7D-.gNRWI
I=1/AaD<caa>6BJeS_B,a?:@/F)C_NXFA^Fe8[c7.G4ND,&E&V@U(7K\TKT<0KEF
1,HB)cWT#?Pa@S2(-OW5A&G__K[FdaIg)6MGUb;U)EWRO-bB/-Nb2)dJI<^5@5:c
2J4E&?6)&&Ld1OI:6Z6@8EfMR=1G@Q96Z2KQ#-GN<&@XWZ2K=T-1S.@T3)+eLeU)
e0bRC./bcHIP07B(LfYB:W:@?[D\cd^2dVega/dbPJO<UTFR3P4<H)3g6MgV40PX
aVL]M94PZV3+4&aXQ/,BJD;F?/.O0Dc+=_(5X/9;.AS\HGHcCOg]U\)GMV9)UFHN
HVCW]-5@]P_[9/=O4<e-c@9>V@_3SZNR47:g3de\V@I>L58RP@7M@>1/XTe,f+9L
-YafXg]WU=-OEb^]9DNV5+.KR7D5]Qb]?^\+.3e11[5;/_D-@@2:f#\dCQ.R7L_,
RN+TEK<T]WD@L<1TKHLg;TIIQ:BWK3,F4DBb6./F>&;CAG0/:+gY+EQ2c].^_eYO
.MRB2bQG-a[?)/J3c4R-LBBFd2#D2/Q[3EB,eO^&cX;K1\=4T[;@UZ75129\:>4\
7H(/L<Y^^4ZU+W1;>W/+IK6\f?&PR38K:b?@9fH2PWN>@bYP2G;)+6UG?OcEL,&3
QM7Xe]L&?Y<(PHa\R>/<2;FLRg:Re0((U>TfS9,=cF^OG.>#ZU):)Kg\L=UZ2gAL
(VTCG7@DBC,+ff1fBc67OQ=f6J53Z?Qe?ZZBVQE5._Z\K,5>E783<;38/+g(/VT:
0Y;&,8KGSIU&[4@P\]L_g[DPI/_1_;9\O>Y-JVJHNVQT@X.H19UCJ(0<AP)d5_F1
X>fVVB3D13VBI9Je?(L>F\bZ1bWHSbOUMDALEVHXGJ3<HQ47./?3-[.DB5@9/PbG
HO)#6D,+(F6F;7U84GK^V?.N#JJS?\@?TKO]SO[P>NfG+55/K<Q;;=WBeXX&T-V?
:AWV@-:/-.=<DG^EEUG=[_e[H<<4/gZ&=+P^L_\Q=,[.:+=f.;A=;d,R6:FNdJ-L
T@?Zd-d9+:@eN-&8e-S69NPZUXYB=#LYZ_#L<,&5NRG2J);HS_5/UI)?/IV.8VF+
H(:fg9JS#355MM,&?W^FfI+4.KJYSQd:;>RFb,UUP>USaG8NL3G>.@P-17BUP8=f
V[bF3&Pd6]DSLUbb_dK0JAc_@e^PX@JgJ]I.KF\=SN#L62e.U(E#P3JT]d_eaJC-
ADC[>EPTUP)bK8J[8;PQ;#8<C7RC[2UMPg#08,00ALIZB@\Q[T>=S^Xa-2feM031
(0fT]O7R1BSS#VdU0R@^^Gd#&:60_,1bXY9[&M]d/)9\5W(WBZ#PbG\(-IZ^80/X
C=,E+M&=<<),,4.8M0a;(b)C1cF9QO3P(1JY]Z_J06&-46FUTaW)JG;^KGVX@.SN
#<JdO2eA=aT?I#?4K9OD:7Y],4-DO7TgI#AUL[3bQ)b=IWTYIP^[eI2R#N0/50+N
dG-0ZHeXC3f7f#T>6Q,6<I<c(^DfB^-1JQSGPC6C<^1)c(&e8c16>EE-(VCad@>H
W)55b6-VKe+;61gO)Qe[X[@@4S6[JSf]FdU359AQT5BW@A]\&LWI0d5N?.LFK4_F
[RH+gSR7O@<UN2;0HT_Y9602b+S+@D,AN8Y@K&;e.3XS]EDXN3b;c;LRNfBF3&V;
>M^9)f=]X5^O6L\SS;bAdZM&R_d^MYN273&345?]3@8DTJ\-575+N?J^#@)1@T2/
AI1_D1DVc@^1^W9H&NUf/9KBI#D:([^8K8R;1^-g:?QJI206A4fMeYa@AJN?YLdU
T-DRf3D/A9dV1:UF=&K>NXP#fH,@Z,2DZ:>M^)9eeR+L[]RXOL8YE]bd68WX,[>=
W&T[LTV+;FD5c[4Q,GPUHdfU(D3bdS=2IV?@;/P6E+#FO5X^#04X,5aHNAMN\2->
,VKO\-?0,A^^2:0\50.>13:ODYLXO>)UC(0]_>GNdL](>W<G+5PbRcYG(5Sg)_]b
622Yb(.@=X?D3D/Y&N+H#/=S/9DZX1G<S,.09KM1Za+4QQAHW?N[0R#]&P>,Ya)2
&&OME?W]XW=bKLJO1P,=5_M:./2FS<O#DWg+>:g(<R-WROSU?W8F6(,C35Z6aYX@
0SQ^^QT@F>^EJ6NVG1c4L9&R,#Rc=9@BVCLLRI<F_[PH72>KZF-Yg2_XKa.>FF5X
a(3.eRZ(2DD39<</5H#R<\J[Td@9#d<IQe;D9,HDb\KC2?3@<4OPQEP\#6T<g;gf
]AJ+;T7cV-a&BP@@7?):1IKeV9KH^ONB(c-a[6OMF/KWCM;EfJ[R6C1e4J)WJM<A
+d0f]#Oac;4>?)L)<U@aZW_^U]UBY(5J3V?Z/U=(^Q3UD?.BNH[PS4]P[<^,JS:=
O\JZ;UXNL19;GcKcRgM]E,ATfg\Y7fWgFE]bFGcd.@A;c@__S<C.[BJSJ&[&YgJ/
;J[d\YAY:7-9eT]G1aI/4.Q]SR^?cKJC@6^9Vb<[&SX99(.JR4>29EAf/Q/C@FV6
\D@19Z>LTeA4JT92d/dd0Xd>cO3_+d1O\gS^E:^OJQ:LMfWIWcVgPYYJdgB=.TR&
R,TA#WGM]FSV=XD+KeK21T3e^&f/,?V#2Tb#ES00V(WQgRJV<dGHJ@G>C3/@TMQ0
YEQ:-4:L[DSF\cfOC-^<J_C2LKDRIVPf,[)8>#?#XP&f00:OC-e#MGLWaPeVb0J<
()b\L=?SK4W6^U+Z[JRIPaP#;dQd2^a9<JJP?D+ZQc#40]F]=O,,4Hc829FK/D^0
3f,MI#fW9I/.4bE>98)@<8Wg&Y\L7Z/.,6bPZWXFHS7W?0^5>GF#VDY37B83-N.(
5^EKN6RHB0BIM)&>NY-S/@8R)J>,H_5dD=I#F;[91@H=d^Ae/M0Oa5LfQONDGI17
CCLX=WUKeGgJ#D8XGJ4ST2WAe;gc9DL^Jdg(IO5geB#/U^7F)adW&7<85X&AL?V^
FBIE^=/aG&FBYCM(-4=9MK.XF<fBHaAa+QMgWTe1>GNS09a@L-?F22WOc,^(?3LV
2J&_Z)&79IRY5>.aTM_LKZ>KXd#_;I0E;SIa00Ig9SF@IW.6_??Y_4FW?\(W-E/3
N.]:G+18FBfCS:eN>]]dWSPS;>[RAAVR96-)IG&ZgJ[GbHJ^1(N^QX]:LH,bgKLc
JGfA<:(cW--L0L,Gec3J(Y9bGQdWWNU,;XRRA62Z>>Q0J^?]QH1-WD;GFT>C7QT]
]D17GX.6f;a,b#aGAQg7.^VT0;4FgZVYf-^OME6FQ^,RLS@MH@+5?8L^)&3M^ACN
(,3IW8L[1Q<3,Z=GMT4a?(Y1f=;2&4^IE2E=#Pf0&;4Vd_RN<7/?PV+bV()2K9]B
R:B?XF#W6GA9O:KG:+V8UXA4^)0QD>.>/1]4Ja&VUZ&8QU/,(fgW6eb#</1b#K4D
63YGg\@KVY/>Wg84>)_0<cBYOW:[J+ebRI:7_8KgRMb2e>.TH-5gWT9OMWHCMe2U
F5I<G\L,][^b=#-NOMT.+SV=86Ga,c^O7Fc-&&JFS2;3_W?:9L<3>Gc0>3dN<0SJ
^8b4:-fQ\OYD&d3N+1-E>>\[R+NOZB7O:S[0E)D3-dBSW=V8>_\0+PXWI]B1-YXA
,N>;WGTS08)6b-<A.(?E)Z@c07G/^7TGVgRVO@:XS14RM49M^f&\cQGEC6_3\R1c
DUI+\g+0C_a:U]CGQ,SeWK,gXM,,O_41cZH/dW=A)c)AGDGUP&daR\@@+J)<\0D0
C^L^-)QV?fT6^C[^3Q5G-fA..AcJVA^.\CRKO5/C@;;4H.3N.2Z<44E]VN#O+0:H
)).SD+^\CFI62&aN3&FWRaE\2;E^.-?]1BITKWP\9R]>KG,9V#FLSFbQ\V.#Pb3#
++;@g)XK6g3O5-,Pf_g#VUaP?BY/Z/KANDGY-^)J4Tg>:LISg+H)\ca@/HER#+YH
.SAFMAQ5<Z:_.;cN?<#<G^OW(GE3^3+&63>G,1NaY;L/F/:g[<8EDF1I1:22#]-=
W5.eOGM:PL)_1?M?R6K78f^bADW>A39A1^NfTa_a]1I\Sd=d(&N@N<)=9>V.D4_7
I^Se.Laea\\,2=F1^/<E(^-<Xg;Ya7d@O6RN<,)>93K>X6>DB]a)F.dN6Ngb>CL1
8A[JaE_+e7F/g70cSgTJEL13f+<gc8B#GM3)(Y9g>N,B&E]Q56+]#aJE72FO>O(G
/7DfF&gfSSg.IJONbN\a_8GE0NN&0/SfYRUg(AGD7DHg^a9(=]=KKNZ1/geb/BYM
(J[Y/>I/>NIO@J[9]a)I3EeC/+ZB?ZCJ8?7L2VZe6dW7A38TAA]]OLb-FKN3;7,/
Ac?Ib1&<Xc_=cA+(:?O\[dP9R_dK,7=R>ROJ92..^^#RL;+.X1J4/dL7&W=#.9.F
TK?^,CL-B^K4CbA@O,E()@c349](@6F;1IQJQgRa2_UTgMd&;\-0CCHObYHCb:-1
;CM3K:H[0?(AEeO)C8?F8NR@5)52)a(g-V^SX6\MEEAM4bTFRH5<K,]C5M(aR)b,
,23Y,,G4ZfbE.Ib;:&W6=OWOLTJRfa[>6X]:F>U7>Z0O]_BVQMLRK(9UdeNM-8A>
DAN-VE494eG(_3:1?6S\fK_)S212CG;Q35T?J)d0(fU:[/A,5F][a8Wc,M=NC_4]
2E\M5#+_fa[:b#BKP[[,_&1MgK5R.J@F&0gaA4NR<6-H5>T]9b8#T62)64PX:F20
8cD#2(U+^0L+WNN2TVfK/+MbJe0Y0&A7-.JR8O[A-CT7]F??11E7??fWQ9M.M<)P
cd/^<1cA4:RU2\5VH0[D&)Q1VLT&R-f,E;NRJ62)=8E9_ZZ+-010=R0S-#]627S5
f]0I[aQV?1c/55+.;S36RE64ZIN?(5Q@SE<N?^#)OgHFOda[JDU)H/NM(SPJY^KK
EM[Ze9Q5GTb]+\&\c3@&;GC1Z7HV/B1ecQ48gfU763,V#]D3E8/4FM>RXQVE1\W-
65Ab@BJ\^:]WE.UW+WdFF#GECF:CTQ&TC(<D4QTQB)]VPIRQg+RJ2QH_WLGYgFWg
O4PM\FT?]P6?AA)T25KT]WN9RNH;3.3/b-eMc0aW]&9A,9L@;@]1>U4c:EB369VH
eVb]X69<@Y..fEI84bC)fGb4SA(JMaPYWYM-MBD@YJUDgFc3cBYH)_6W?7U_dd.0
+d43QOCTZHMTNAb-,P[ddEDGe:T?S1TNQ99P4NQ45gAP<aQYPR,]?[/AgdLeZ[MJ
AB.JM5R38NSRe^G3AYcAA,1,21R):&D_agVRWIe5Kf?Y@>(S>W#MbDeDQ1&_E2@b
AV(6<D\N=S6J^:OR6-/05Y+V<7@4&?YD\JW?LM(9N_P/P;UaD^45cSaM^>A#Y9Tc
.5R9_C^[5K-&?/]-\1(<C_SeF.-YCD+0bLIR-HVg=5@H/KD_<;9I[4K&\-O;aBU-
7L0GRb]AYTFS,7^48I=&KW45g8ROVY\7US#&dSOF\XI2^:@KHP2N^D4TD.b9HDIA
PIad<CB_[ZH[Q46XH7PP1<I6gN21<^IBE)TS,4e<](5_a_ZaUN4dZ,Z2QU3O(ccC
4&R?ATPH--HKa3Z6:FVb.fQ@8D;+>c2Z?8?e06CK],AGI4EJ^DV5Z4PJRf^C9(;/
WEb)?05QaVFb8)=_)faA1JM?O3)&[>:R7c0\Vd5e3>c[VI+WXc5fH:E_4+V,N[Ff
N,1@^OILN)AW,g:N9ea8XH\/DNJ]I1?IdPWIP^)c.:aVH1)SEDPO..fdP#9A06=H
IG?_f+&RU7LV0WE,e7Y@NC(IPWc)T[?<JbBWfaW_J#89[AW#HHD)9?)5:D9ScGK.
/,,,_LW;I.3K;1OeKFUfU)VSGfb+b.AZ].De6(Q=K2eAb]0\OLFAPbF32K6]M#]N
M.74I^&HR;WJ)J\X1,X8^E8fS[+FJ2Q:2_;+QH0<WAf&,H4<5M#-T/>#,/MUbA-,
P<EH]7+a0Y\8b]@0@D,Z9DHB,TU?5>60c83ADVb8,2,3.QT7JA(1Ef23/PTW0C5\
\^;?;K+d:dL=TEL(K;1f+5GSbA,F>QD)@_=P<cafF8RO1O^,&[J_2BQ0^/&U7Va4
9T^\4U@:#5^2+@X3C7A&QR<:I<8LA]D^71X)?\B7f<#a<A8bCgaOQ_V@P[I+7,_-
/@]#M84@8#6K>WaX>SfUBS[J;=;GN77MSR/g-?+;K9ICKRO.7&U[4e#dG)T:PIKD
cC0YNK@8gEPLG6\cC.R5@1LV8M6WGTffQ?U=2-:937P]NH_--3X8&9QH-d1YTCX[
HTN7AVT=0AL?7T/CV<6EN_M=QS/f\U\84^-D+fAJY[Ca&a8eZb>d9dBZBS=f>2GJ
NO,(TbXA,6\;0VFPF;&[\8PaL\4b(B6ZN-V4&WB&.^&QdC#Y8cUMfDJ;K##MgH?c
@6@A_KeeA\4d1&Y^&8HT;WKJN;\6d/>B7II^?GYQ3e)LDaK5C\&g?HD_gfK#?SaJ
c>F1H2_6;CJ,\_gKI;&.f(d_.HaI)BY?=R)UacJ(&3-&I\N84XNZP1LYJ7fUHR:>
86TB8@6K)\X@eV2RMW,DV,Ee>TZ4.B3Eb<J>+X\V_652[>4O<1RLf(>H4e2GfB\A
2F8CLcc&cIfZ&_e77Sgd3KL)X21eYd:7gZUQAaK+b2;2ERf:ALRX39KT;AM)\9cN
\XK+gKaa^bD-bIY]7DKNH2>&HKY^(Q0+JVWHK#E5HI8]F6)1WFV-PMAZJ56RQ1&0
50)d0T)<CD4A:gIW45YfMc>)O,1c.DPf9XC+,EU1FP29eJFaMJXIF.IN[d+L7.C[
;[?16=a6H)aO30=RgXY]RbBAMDbN+Y/.@>W92/T^Ye\AWf;faI,U2#?#VEOLNR9A
C;6I(-7]Y@4\L6?4XNe7PVKWLAKK&IV@UEVO.4KE5W>>^UOc\;Pd<:8.Xb4f3eD/
;Ga)VJV^>IH5D3gQZ#LFK3+Y/@9U:2c\A#cM1BG;5;UK[eAcW6N,f\6WSfNOd+2I
NZ/4FeSA-3ePgPLJKYbH(P[B8,V(/d9N\Z\VZ]G]YD^+<?+XF#]RL0],D;GQK:Y4
4OOHWMIL7WfFdL1,-Wd8J7=6JZ+H6JE^I:VH47Ya^4CT/J];&2d+]V)<G4F.CQ2/
3#J)W4NBcEeZDKA-U&QCGb7GBV&a7/>XNUaQ)OC1OaA,4/A61<ODY_-ALM,.<SP\
)K=[P.E]X6AIK^.3-CF85JQUa1#4,6<AD22U;=8&8R4H8[WGgcU?[0..EVUbd.7Y
SH9Z&:YF1065>H^,<e14;ffQ=c.gf3(./Pd5,8bB@<8/82d+dNMTbWe1;@ERPb=.
-GI7ISIB3@e,eY+CT:Z6/740C(64R?\649<\TM4eV9gF807AMPRV2YACU,3;5\2N
,TdF#^daFc#1a44(\c>XXf^E4RPY[F1dd,HX7-cZb4+7Q4N>K,.B4HR6[RFDN:Y3
2(/U1@DEH/e9KZ9VZ-Z=YeEX\->e;>B9IIf4K:@MH;EKXJF&/WYO7CKZ_b]/].=?
c96^OMgZG[PJX64<CcOPgU=^Fb_6V>FB+0eND[O4#c2ACC^>XfX5aP@gB4f_8F_[
AZ6_AHB,fI_YPE,_.YJPdQ>O2YYD]dU>CS3JNJPI9UG^KL&(PD/U=2;IYN\QXGYT
^M\Idgc.ANO+]Ia7gT5<#V6cYa6^V3GKWEMG^JdU(72.<ZH[=[(D:[,\8eYOT0=9
.?VJ;;13@W1IUedGTbKBLUc^\W-M\#C)SVCdF8).6IfKO>.<+]@??1bT=f@^P;EL
A4I0C/\cX>CD-9D[5=37^LIB:C.7VaOEQPM15.5UR2+1e4G05ed(2PUHRUW8]OKe
#L4W;aLe()?[A6^]Z</;5eTL6]5C<)cSL:)SJ,^FTT30/_<=/d^/5OgM\)F^DB&f
NH;3(e=.N]@YF]3HbPE9+JZ_D:OJ\V/HD-daBd#V_5B>T1T;+7-9=d\FDaN#^UDN
b)5-Y\X,XSCWL-^9b]TPgU(F3UbB.a^0#S^9aD#1->E>2LYZA):WFFF&OQ69?Jf:
2X^RcXQNc\K5K#.9gO2JY79_AgUN1-]MI-;3dG1BL/VG0]WY0fD#H=]#FgQK,.TI
2d8_E>AdBW.f,0SHDN@<3I^A[(V:U[<RPLYZ+=Xg_P5EV0TN@bcMM[<ZYEDg11e,
VVUH37P=28I3^ZB2fH_RQ(@?BPVI4+f+:)Z-^E[IZDCeUY[,TSBK8]:4-2+FYXdL
b1b/Ng,WT+5<d4BMb^?KL_/3a;RTJY61^HbJBI7-64fZ?5R:F9&Z&]f:.IK(WXgC
A.MAUbUOc6^]ae^-gU/e+?/Y0A7CXUL>>S(K3L@E#7]_\>7?2&KbBOAe]Fg2A:1R
I/HfFQbfCFPGbF<B(/<MV]P;WQ?^aV?:&@#^K</egG#9D;IW&+/W)<3?M>_)gD-K
++0Nf(F&&]^O3ZF.U>(WceWXUD_AO#CS=ZU[^.5#9QAX&KX[W=Z#RMY2NS(@LOSH
[7bGEW,732@,NUCMZEG:(Pc5(4b)4QHNWXaUegKBFcgaFR+TAPT=b]H&b3G(dE01
(+5F=J@<:R+?C1UZ?Lb?TE\SX2c.gFd?8J,I>^Z/1F]5f3^f((UW>OF?IaCc]f_g
g7c8HV]\C[E]6Mf^.Z[NDbSN6P7C/X2838A8W/^OP>G+(^VJ#UYU<#.I\d:)\Te(
6R#e;:gI5(9+LUb-X[QF@U&JQD0I\BC/2E.JI2#/WKfd+I@LAdDR(^^IY;\WP^<e
6LV8ZMc]:-gGb8?[F6A_JXY?=[HWa4ADDgW3\Ncc8XV>0\bD3S2H:Q[-CdeYQPBR
J9_JWS+.d?Y798fPWV2cPY[1)TJeTWMJ5ADc[7HQ:\7dD=4@B[LSBJV_3E&9BcMD
Kb/&gG.,<;QNdR>4,QTWSMDCGe18>^,@1?]2WFE.1WbE;a\6T8RK5c(dF98.-?-6
f.5)TEV<8DPN@(=1;4<V1#4e4FaZB)[UBa<=EU3aA3cUFWgO9:.>D-AAWBTDO7g/
,c@=&;Ff505g=NZAg>Ca8V?^Ng<P+]Ib@IBX,UB<GB9\Y_1)8T/Tbe^Ib8.I9aZ4
eEdOObAOH=IfgB=S#4d=/VD7,KS/Ye>c_:M=Y)180TH2,3DR_XXB+J<ETNc#7@XX
E\U0Zgb02O@RFVcYRPP9KYgD=<41WX4&PPfW/EHP2b#Q[fL/\C7ZG+;I&X>/2SJc
4M&#LN4?T,2Z=],<R@88_@XV7@N]\XK@bb-+DQ^LB@YfK931TRLALTf<@Uec?b[a
I+B.,g_(NB6<Ha-Qa:87C=g4V]<6E6^)Z,M9G?c6J>LHcXZ2cHJ&E35ZJY5T/6]C
RV<)B>fB_5(_?FbP1JSVYICY72/#:CGV(#[F@9XO>#OT].^Z]NK+/VHK\YWM8603
<RRN30OQBA7>?XcT3eG1W(MU<T^^+aeSDWVY/7JL30Y&4E)[91\3f-BAAJ/TZL4:
X8(&SSMUN<)EaL;L+.&M6eX<NSbc)JDb)KNYU&4E]@K]1>EadfJ/FCBAK$
`endprotected
endmodule

