//############################################################################
//++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
//   (C) Copyright Laboratory System Integration and Silicon Implementation
//   All Right Reserved
//++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
//
//   2024 ICLAB Spring Course
//   Lab11      : SNN
//   Author     : ZONG-RUI CAO
//   File       : PATTERN.v (w/ CG, cg_en = 0)
//                
//++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
//
//   DESCRIPTION: 2024 Spring IC Lab / Exercise Lab11 / SNN
//   Release version : v1.0 (Release Date: May-2024)
//
//++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
//############################################################################
`define CYCLE_TIME   15
`define MAX_CYCLE  1000
`define SEED       2024
`define CG_EN         0
`define DEBUG         0

`ifdef RTL
	`define PAT_NUM    	5000
`elsif GATE
	`define PAT_NUM    	100
`endif

module PATTERN
`protected
ZLH^[UT\41g&E@9OS8\B0[HeEa3(\;W\DV[fU/A>JUg5_T)B9SRb6)ebY@5WR[g6
JfOHNW.H9PH,fQAS1[(/V?HY4YR7V6S5\.BUba[I=E?V;8gE>]_8IO-7Dba46EAK
_[C)KV)GN8(K<^AKN@PN=>eA)17-U.EOI5=^]R_<@#YAQF:Z)=I7B(b.MMQO;Ddd
PACW7)8cK]RQ1b9U@__[T\f:&M;Xa\H4BT+:KW910&N:=7;f8+M0+a_:B59fA4S[
IcL,?(]fJe;dKS[[)^E\N&f6JTg;UB_0GZEb&]?dZHbMPVf4L5+9d4;K8d@7-2,-
M>eE^:G[<([RE6_WKBQ10N7:]X^MKAd+6I\b&E5ZAaOY6HWReC3/Z)PVC[0e0[=G
W/@1MGN@S2eTUT(7KHKaUHNe..T<b?g2RI8]Z+XX>-g^P5;Sg8Dba(R>\/F36U1Y
^8VIC/O/8]GK_e_gXgWPC3UFB]A9P@#DC[ZX^dISS,\=G;JU3UDFNN95OY2(M#WS
?Y5:OZGOa+HMcO8E1/;EQE+RFK@JBU>&7QGZCJ=g0V#)DQ:<VD5QPX\=XY@bG,(F
]YC\>2c7)/2FD_EaPc(_RN);:WM6,g:>KIJCXdZ)Q-=5b1NCZ4L#<==8M,+&=2@-
^NM>C9abCgM#-1dM;4gMQ+Z8O3\c:Yb5@[\\3e:.,aECCR4TPKY,gAEB?I4O>6^1
M=>)2-#=bLFIHGHgAfJ(>DWAE07DQVYJf4T06JO>IT567S/Z+Ia-GYgQH_=WUPY&
V.JP.Q.EgB(O]X+JXF)Lc.S[^[N>\a?d<K)_1CQc\@[J.OK]T]Y6A=)2c_XX04OQ
c<Q];_?)Q_;_=^,Ff98-3C^2EMKHD=,1AdOa>/\E^&X?9VFLVG+C(eJF1)Kd.LPY
A]cEb:cc[B)XgA3]]OCDcaS<;G-Y,ZP/G59^T^[#c,K01_TD60<R(60/<dGMF0.?
CDWdJ0?cW[#0@ETAR-7SG\g7dPc:ZRbb\#.H]KKbFBT?]0):MbG8S:?UWN,N3WL/
51GAS(,M=IVac+E+d@O^([Kb9&:3DZfMaPKg>-f]?DbGeKA7#,]7.317KB0/;/&P
HcEHHYH]934B5NW&@]0/\\AX6)?be^(a-R&MC42NFHbB4B)+N/cf]YLJXXN4\^V,
Z:X\KD^eAFbJB,F^&#MG9.GA(OG9PO(a3+3\U64bM^]A8=W3?-UeKZY@R7e=\7b)
gG?4?3JF+^7ISg]:K0Q<54JYQG@fH_gXA8MN[6MH>@)<bcaa)\^I^3Ba1FD2,(<U
WDR+7<Y/XI5V25D0E9eN8PSW<?_KdP:ML1/E+CYBGG2decf<L^N5QAMP/^0)99U6
2=JT?F&1\fg;4-dN49GM#.JCDfQ7UV)2K.CObA<#U(WBOe>UAJ:I\c,VZ_H:d-#c
.YG7T#@4=Of=52B+OZ<9gfUUA2.3X??:<VaI&=5a&C/RFF^NMEKQ/Yf)cWDNLX;[
[gH^FJ@D4=GY2UdPB,AdJ@DKNA_84.:W4^6BgFU=3aNL.g/VX[1(SQ1SaE#R5eTG
69TbZc[0>--DY<Ya:aU@P^Z7:-Y3ZRB&L@C8J?TQ8:1XJ:>2\[O/3]4TDeKgfa^a
9WH3)KB1/9fHP^8.05OA[6O=T/e/\<ND+)6K:]fC9VVX?>GgJ7]<R#=P=@JBAf_b
UX;G4TUR3F3a#]0QK_A\ggTI5L^+-6A>52(67/V>L]\RXS?@=9B(#?e;Cce8M99L
Q)Sac<3T6@4XN^7fLB.G&ZP1gcG@1=_KB=PS<Y#O9H7e4Pa0-]2OOCVXGW.Tc-6V
+6<K)cf(H<T#IfM<?[BO[AQ;N(FQgePTH#3HDB7-?O3D[QR=5@:4DJMMMMbHc,,b
?]CeH\8[]dC(J@2>:_bL1H(@eCc7de6.6c=1SA=\9K57T/DC,BZRU@)Tc=e[>P9Q
)V0S[<J+Kf33=/51&gg7DDa5[3?CYH(P7RY0Q.JUQ.dg8gF/f3)YEBCdBA,Le^8W
TEI&FIZSTc5/GNT#\D<-99W\+aO4g^aEE#Yc^X3b@6DI]^2130OBT<e.S7)>1M4I
.?9,ZHf0//^[_RSQf9RU22].ZF2ER1?;UPD2]2c.3G\8,a[[(Cc),JJ?QQC<,2O]
ELTX<c,f^_d2]FPQ>WAKaf8\S,&0E/bV8OCNbNcK3QgBc62]eJB<AEeQOS-MGb<Q
8,KG[SE;YK(U8B,AR)Oa3>+/SUBA+@E0-T.<35A[5UV]>KKS+Q0N8^VcC[TIf,U?
N;YffO4XAIN7>=QSQ6Kd/Y]0dN/ZPI2&N7c))^ffA]XLc/]1&64@?I6E+6<8AG[+
F]c+Q,T).6NJ5#(>Y-L>G9ME_JTb//RfG/6PgC-0&+:86A?L;Z#;eB7(YBGbNIec
\09TO^?G2Vab8dF,-#POecY+PW5D_+X_b/&P,H4G\HB1K0D[R<cM2EI3E&NRYW=3
9,e2dZY)><R0)dDe+66AC:W/P,/,f[.f0M_=TQM,EDa?;2[EC2HLPM/Q.[Jb5MLG
MMa,P#?)+1KB]gdA[&Ac60Ze[A3J:;M/LK:OXK8P1FV]_:#L5,Fe>c:[9#)EZJ(N
PTOW+[TDRTPa]b007[H_0+5@)dGAYK\>Y&@X3MYRSKNK)XJB)fc6#c/X&7^(].O2
;U;XL+T:0H4QU_4@Q_g9&YTH4T0<K+R);DOL^6+(A7cM52/Y+_OQ0^T#]=D5HU0Y
gMH@@#WO5P0O6OgT<e#QX6,eF4gH.];I^.^KY<KC3ZO><]2EI2fdVER#7(@1EBL)
-ad@CG#(?QRJ0[2Xbd];[DAdTF=:V/F^-;Ze^O;Q)\D=D@c46WUPa<ZW;f\<Z6E1
^-YN?M>2T\>>Ca.B&]]Rf&6Y_,T,bbP[,9Y&\0fWOA16P?\9GTXLad30,YZM+OI;
,EX<=/9J)2/_5CF;6OX\AD8#,e4gYW;,&8.&][2b6OQ:^9dP)V?g@VNR4KFQZBQg
[e-04#]GO?Z)@0\^F2P7BW[a6H;-S^7S64OD?dH_]ac@C/cRASTK+U-@A-dJ1>L\
g[#P\4\--b_(;:94Ac6+=\U8eGag&AfQPBdU-9,,S;_B0@KLcAbAb01>Q]Y5Z=P;
+B,]Z(LPb;,OI[e1Gb,8L0=(/\#<27>4eZ[2ZF1_L5KMe./ZI#L/O#+e]O]EU.5+
c3P7^9T/S23N)3O&>@HD)Ibc&^]PE_1JeLM/g?^DPM.V-346^@@V#>0U/fIRB?dH
3AHYL&e+3<.8+<[Z@7g?T@.PKL2;7K5TIW[H?ZJ-WMAP)C&f_K)VcP2&/a#=Od9G
c4d2+Z/2MFC8eEe^-fAU,.\CFg5AgVf,OS^RaBZ/4(XV/,:S4]e9/f2/3-?8DAVH
Q.WAT39&-?XW9)g@N45EdE88c,U>SgAM(XgMUP[baU0UPTPY-Y.TH,fBWfdMc<U=
d/C0=N=LB<IH4<F@V?=(0/E)F;_^D&?@bZa9UF3_D]UcP:^OcC^JRQZ07CAQ6D<[
cB\)).CFe?NWRdBJa8<E;O]PZ7TJU&LV@Q16:#]c[_0L+P2KF[:fP#L;VLWc9X=B
>&eY4U1fJ01?V/=(/C8HA>TE9T8Z4Od/dT&X#.?^=0)-f]H>YYC^PR5gf3(RZ;O/
)5KNHMI?_BDY9[g_?g22+f^gBXGL\]M\3b\ge)0=SAU?@BJ&dbbWc2L:B6U].A2B
M>[:R(,gAW7_>FLY_1@Q0AHFS[U]8[b@SIV4<LT_N/;1HbK0)K3dgI77DHOTOW<F
b9eU&)3K/&7YEVL(U2=T&@IABBVaU8WT#W7S),ebL4SYED-RHM<48JT>T@L6#0X\
9.4]BE?,54bgF<Y-K\48SVK7Z_7E3N9,e\>Ie,Oef=0g88M=UL:Xg]/9J8BA#)3Y
CD-[Y<65aX4EUJ[NCPd)=Ad5<.O[5_M[Cc+/ZdX?:WO6A#QJ6Gg]g2Zb2.YY/I,&
g6V^IV>P7XLA\28A(&Kd=Ig:8dGc[_-&Q#;>e)G:\+@0\:>R6T.OVZ&@A^aSZY<I
>?IXQgIc9dQe-MfGXJ7)JP.B>A)0_U,:B8=/VGLG>S?/;Y_A8BCEf##OG(75=#\b
CEe>=L+A;YJ=HUE1;Y.AVZg\d).;(Ne4.[FDI.0).M+@c@BE4=<-cQ2eEfdWR<]<
g,_ZZ;@1^a\<aR-<U,\JT45J+#:94JTf3&#5&9B^cTN#J6<A]e^;?^,:c6/^=SY3
J2Ug_V3M[>f;f3,-V,2TC#-\WD[?=I]@RGF/P9OYfb&]gNYcV(7^Z/L)4MJG5TA7
1LWSF94CRAS30;T^f#]:C5ZQM#T=cTgN5IS#?^Q?CJ<[FIfT#+TaE9^--geb:O->
D6>9Sb(X8)#fSXW?(A;GLN+<8A?<>0_A6O\;W4CDZ0@9a;4^aZ7B.+c+-@J(/\.S
7M-84BUSPa;BSbg,;XQ)g,G6>&.C[c].<BbdLB)=Q[])A2DE#C[0gIe&)&FEENN4
7T\]OVBF/A855IL,T0:>XISES&B+VLD;_1=47W\>IPF5IE;4Ia;L:BY<bTCN7R^O
T^(>.0RK;W6<VLEJ+&=d]^Z5bV72.UWH\AL=4K87Y<C23LZ./ICX+;8SQ7,F/ag&
AWH(2.VG&2CW[_/=M>e;S1XYFKT.-3R0W:F+WF?aeL_LX(bQJ,RRES)E-ZWV(^ga
,M26RLd]?XH8404,A1V^+K/F5>7<aKPGeCH9#)5\=#)SKR2\@K?Va(b8V/H,D#e^
Y_T>B0_CU;X+MUfZI#<EW0X>d&<8-RBWEB?;/B.^(7(ECO=U#4::aKE&W9.F4.GM
#FF-[=(#N&J0,).[?.@VSNcRN[5#]#20RPO0?JSMZHR.)/_^5<Ge304?/^RSZUQ4
<=R=+I&:)E#FY<R6<U#bfP\WCIRG)&d4cD<B#QV4b1F1dT,1&KPR>/dOBQ.O+68@
+[bgdSDZ;R#_B(PR)@Z21/F-BW)N7fcM_Ne1eR7UFIBYf7egUH0Y9S434K\Q]9eA
W&]=XRW^N_836O^\BZY;T3Y2VS7SY+H+.4]TXR@+]QE@@1F5<LBeS6U@M]4DK=(P
JEUB3R6&(Ld./EYNc6c@D4ZNfWIeNT_NAY]GQ4Hdd8:bW?D5V0eYD\.T0C#MK,b0
T_,ae>9@3WQaY.<HLQT?F[)I@88a>)8Dg40:ZAT^1VO[@W1ZcYbc,9]7S&^+_2>b
LRCd_Y2e>\/:6#J6#/JN7E1DMGV9J(A/0LX62IX<KY.[0QOg?7(:HQ#DCS=+2^YO
Q9=IE54\>KBIL/IM65Z]+]T.F3<^0P#c=6WB\\LL+KV1eEZcWWVLf(ceW<(-E?Rg
-0;&-#S+cfWd_bB@3G/?PB?4-]OX>^Oec-<[d=>4MDMEHU?C<UUadK-CE<a[XZQ_
(Y?8;N/Wg,CP;UQ\RSf[B#>6TC_MBE&5PWg,7EaF,:a]>>(30?JZG8VNeUbKSS32
4g\IT:J[3W@<(8QdFdGc;G[L&F1]8gfZ74[]#9YM33029/]/]YLO:^g_]<2W)eC]
R(BXYS[_BB2@eI(Tc?V)#;f86M6@Z7UMCe03d3OOgXOZYAF.MR9(=Ma#(-R&ZBQT
Xe\91(?-(LbW&ZI)H=dHCb\:_QAL2ZEPZ+36UEa,OH7KVG0TUJFH<(.)JSI__Db;
/E;bGd;QC0QE=NDR(_c;ALe4Y7FI_\X99@#<IQ&T=/LEMF)BI,7@K8=Re31(N5.O
X6Af^B8JJ>@</SJ3f,@<2OR=,.:R2J7bT_OMZ:D.RXHe=3)GBcGUKa)&&=D#QRYe
d_[_B.Y-FTZ9b45-568)\SdI;+6)R:L)>D4eFSdLL@dg<PXN0e.9-EAVSbYMDa:(
#cQ]f5c<)GRNeV]1eeK=#I@D1?:EA;Y0/eTD@TZ&\H#E>]cJR-K<&>)/C??+=L6E
;__0G0C/68S#F.G+VGC_GO-]2YX6^V0:49C6CRU=#SU#AHeI.7M0+>8dEGXeRYB9
&][47P[#+F^1A98;?=]4L2XE;]+].0(3K^.K?YSbW:64/eQ&/DP,f1(6g68237Y+
OLCgL)W(Z\\U0(&/&4L\94Gf=I9Q[S_?48@0),2Z#R6;9bAG^2bVMRc2X-B8[O/)
=KW15,@?).d4g&TN-?:b[0]X\)FE0^\J+UEMYLMC\^S?)f6bL^FMV_RE:X)T63)?
K:g&@:TT>6)M1RS.8-L7e1DID&A90c\(Y(K^ML&@5_:N:#Z2_W)7d_.Neg#Se7f/
c0U=XR(Tc^Mg-K4F2__=./<)AY9=Dg<Z70/VCLHEbI+SCaG85G,/J_f)>NKA2Y0M
Q:OM2I/-I=eGWV&8)B/M>J8=1@Z@<8LZIP]M/Eab0aERK#LfHB4@STP:4TI>O(gN
GP+-AgI;W?]U6bC3RZ^1;HY<H#a:E0c\4ZP_/3JKI-A)R<K+4bO3N<MgQ33/B@Q5
I4NE^\=8V2<&bbPLg.EF-(F,-JZ,[]PP6c[6FG\,c2((J96U?Z:b\W/]W3]=.5bM
N.PeO5:U?1G68,G?=f,5f7VQ6E7X=B\D/GdB]/FJY0F54-5KP3^1PR-Zf3UDU>M#
#)<#4(LYZSISH_S30GX>#H\PDS=gM5\Nd9=46LT8D+ecQNeLbO=HE;DI8;N/P5PP
=6);6KX5g@K\@?d=6f-,XSB9DW[DAH)G5Q=+_4B<MNR&JBF+e<WSD1G6gVBb<5]L
[?=^_4C1^HZBZ?\,[BS1Y)&3A>SIYXKJ#QJSDd_Ra\Q9>]WgNJ3W#>9cCQ@<M#W(
P9EDd[A)BH68S#)0;LG8D@?fF&+#4@X&T.UL.TJD)OR6&?]QOYBY6.+Z/9(?UB:[
[_/W::4fg;19&MZ4\<=];4Q8W.VLVYf^GWSTEdg2aCg[MYcGFeg1OU\^KB/?+WQF
UA-_?R0G8>22KcRAWX&&/MRdM@2>NCOM#]?;9OT)WG7Z6Y.1V#.6WR>U70_VB>KH
aA<ABQW#J(^6V7F02@WKV;L^[6/;DTDgb8?Y,\1L]_H]PI).CFTOI7627VfWdEd#
&S530f@;#OY79^IYN0;++,^<f5JPCK3G:;(O\2S=U6M]J&PQ[VVF&fT^FHGAS#OZ
1a,KB(RAbA30<V-]=#ZK4SW1;UHFBCM:QZ8^.W&SB&20aM4@RgMKZ_2e:W7SITd@
=Jb)((._D9-MaP6Z=M,U-4D^e.O8JPBcW5#7O)/H7B)IaMGQ61CTGSCEgDCX9X>B
f+83fP/V?N)\TVWA^=\+:X>Wc4[P-V:7@Y)NA)d#-afIUfZfdZ]/2E(2Z>F/\g_2
:U4eW_B0-8KHYFGVGMBRMFA(VZ3]4b0SVEUG>a)/B&(/g3\]IHC]HM^9<J-D-5/4
(d,C\(V?[.[DRGegVO0>58[19g[95RB^<O/D96(Yg50Y,fP#X8<M,eaXEW9;Z-K>
PA\L)B8N-RHQN9KLCUOHML=5ES4Qd1dMeJACZ8(5eeRZ.ZYb@>-d4XZ@FOR#FSGO
HfbJ\+\]dF-a>8N3a;X5H+0S(4a+=;O\\cR5L:3&GP:XG8cfBAM&.E_<[^/OZE9&
RKIggT40@WOg-5W.(;G@<H\@PO45S7W[<.?&=#ZC3KUbPVK0b77?=+XcTB1^:X)C
c@FC;S.&N3?T^-bE<7(Xf4]S+V3V5<FG)<(#eZ/g8E7J@7eQZGN/dgdMRUV-La6I
+S4\Pd#DK1&A)Z:RKDbIZ+ga;1RK.0L8.FCABHRJ5dF^)e_2DOe:ANFK].[#FO84
@Mc7B:FI@);<30Ydc)b;cE,1C0>Q3-/U\#1)Q^U53)Ta2V2H5K,6(]=T49O2U9]/
;I(9e+0X:O\9\ZbM^VcVgU]Faga5?8;gcNH2XQ#5)LG[3&H1fH#VBCV>VPX8[33L
XJVCU[;0\QaK0Y078]#HK,I,Cb@b<BYe+fRG.P0eLbX[fTRXZbH#26SZ,9CBG>eG
F>8>;2[G8.A6&A@MJ1]A?9(..Z;3c?--K0FD1=d^E7a=Ce9f,,Dg_^#7O1Te\MY=
V;W&4;>KO=d6eZCZUQE-A0?S&67U]PM:Xc[+YHfN9Ig>#^:45DGAREa(WD+J&1e+
^Z7/a4d,I&?c-d;&P39D-KAESL&U&(f5S#YYUFbS?9=X?f(]-7:0C(YeFW@2]:>P
gWD84R?33?.DdDe#^80>XdG>b2deU9&a(fcLNIg0Vb#2A;=)@b@D#,e2:8Hf]JDC
GbJd0fBgR@fE[BS2dZB#a]VB9Xc2/(Q?D+[>:-=C2)fZNEGY/J&MZQD&(adf[^=Y
:5@MGNSQcHP\DD2_Gf95I.<A5S0](A,4SU7d1gc&4aQeAGDc>ZTQECK:F<LSf5E7
T;J6ZSb8_>5CO/FRV@#^A]MH9-U&e?XC?+X,f]/OAGL5EOY58:SeBRRQ:,.gD2H0
W1[cKKNOM<]e=;WCYa3)29^<b?Gg#O_TFLBL(Cb^Xd@c9J3=Y88C#L//NF;]WAc0
H[-\)7_MF\RJF1O:C\0_@9aZ4W_8L#^S,&9-+Xa&^<OP_57_HFRC3a)<6PM;\R8f
X@X_0/LKKK58,6^GfHH?[B69dQ/H0<_aSBa9-O)b8e/@5S4\GZ9MIE_bU,+YeC>F
.OWII9GV9;YO;.9a?/<X=_Z1DT=Jb0T/P3T4F,:QGG2UgDSTQL-+[HI=W8+;Nd6)
gH8S1aQBU/M79d>>RS4).@0?[c,Y8=@E8=?,TR_H@4<IW#[(f/ORbH9eK5S6ZU1/
:-JbIEQZ;f+K+PMgE,1YJ?+?CAD8IR5/1,4AIJ&dO[59.2JW?5Y#L6<0@W[(97L5
/7gaMTg3D^EQL/ACBg,,Z<Y/D0\^eQe(HG2P&)3H9QU(cTNUO]B2J_26.ZKCEaS(
9.;\K?Q\bW163OBZQ6-4WJdZg,F4E@<RKF.N=T#JLd;AG[<2HJSD::J)TUSQ\Y30
.ZcUfRT,B,^FIZW.TY<0;0V31.7O\O=,LIM34Fbf(P_4H?\0Q/-WZfH&#ST==@.>
ZR9?\Ze:IO.1QED@R&3MU,N>R,1:e(XQaB3)N9/6R^N^^;Z-Xg/0[9#37?(2Z93-
^gZS84JQ,Ng],L5,g<b?)5Yc7LaMW[?9b&6-I+QWT(=QUbG7>))a#-O>:JM<J>WC
Gg/]N3G@Cee-ee=.BN+N@:B>RX5?+2A:KE8LYL1@I\BYM&B7944Agg06SUNe9#<+
;CUR)(4D7+UYW=KdG291A2+3aWe@R5<Y0P4+E=X9<92QU1F&MX?B>-Md_\a4X6MR
I3(AT0=:e4K\7CB.DF=5((^7A4FXF&/6I,\3X;5Z(J<_We9W1UCFPTS.TC\P900?
HT6UZAQ,4FNae[3F6?548G&4dQ0W&KX>SI<d#?DgV>?<Pe?Xf<IKK\MN.Mb-g)UR
@2b@^OJ7@-+PAO8CDQ2d^.,4F/4LPPMXAM_4NV?:Rd-^]S5+A).,aaI[.=L?V8,9
UU^/f[W@.Q/5b\M:)[Q/FGZB,>)Vd<L^Y0c&DDYM8(NGL90B:\Y\CW[SP8L8f=\.
=C5I-G)&<.;1[[]B5Q?F.^/47J,H.>)IZWW2,YA,1F(>1[_;,MN=[P]V?:8cHQ>\
^QB)]gY,\gIcN41G^.]MNB&=;OSZVD6fQ\++QHM;bS9L6IPF4@O(UB,@E^6V]RP]
RQg=#C?-=^UfY&[&VQD21efA=)b.<P/2=K>C1Gf1>]GU:K-W+M[bK>4?8WH;F++T
9=NV4S.FWCRSTHRa^G]OfJc&ZDNVZ^OPMR]TM[B1VDS2M?X/4>TOe.ZNc^FT7(&/
E.M.0SfO./ZQ;SF\1;VT1.WL/#D.Y9O,7;Q8UO6&TO>ITU&KY(;L[C<D_&B(/3[e
/L;c._dTDW[W1A.?L8#b1fI&+ST:/A<EEfM8JVI-6N5#eg(O:)-cXd>V3;HOZPL9
D.)]9I=G3R8EM&EF[<Q\eKVL7=I-ECC82cZ>1&cYY;J2\d##42EdLBcc8&fX3RV<
BH9d7f4F3-#4L1RCZLHB=S]LD?0?cZ>VTg#V(>fW=81CA=Z9Sg&ZTIV)f@-5=+^Q
O.KRUU-Y8aR@M:X-WQO_F=;^]5dVDf3#PAe<C^HXEf9JW&9Q3#F+5TRUGI1XB5Ja
X,6RD>BZ&9(fdG4acb>,_ZRB7\:]]U6/c3>-E(]#N)b6)+B+b[R7V/Y>?0ZSf@CB
;65_:,Y_=I?H(EGU@18ZX@WfQ^J8(-1;Y\(-YX/84MT\[6Zc1_S@(Zc\HRFK_TG@
660[H3BO\L>=RWUK&A8DD7cE+8NaR+\\E.WW1:TS=;YFM@Y#,.;<faMF(JgO>EPC
La[b/;P#Q.<gO]5,I^T?00?ge-[07RB)A0Y0;&:Z1-]94caQbX_[X).:0<H43F]1
=cHBHU2]ZIFVPW\=J>A7;b(=C,Q_bFB2#OQ[Vd_ODXBJW<?-PYfC.MG&G5dT2G^C
GOIM\//D,4]8U0WDV2E;G[A58.2dY6V4+aWN\f<],S-5I#(9]@8#9:8,bEGTgfV@
?W.7Fd>=26Fc3XM2+AD1c8Wd9_Q?CCbOAf>NSBS=?_<.X>Vf.eE5F565[SXcY^L3
gMABe#?1[./LPJ/U<@[&B40/5fZ(RbVb#02;bdNB,H2P>I_Ad52PeYEH-=7d;-6#
/0C==@,d/ZXEG:_R=<41\;BcQ@0[aNK]=C:;MD>1N>)#:,Zba8=;b^TWA>#=fNgA
5V9F:QL:2@IN;bI91X=1RHMg^-;/beBY21FI3E:-U-AUC^&J+H<R7+@JQd9d:NeW
2L@VC^fA42LMOO(aN[\9:Ga,(=8&I-eYXS,gVUER1A:a_ZKI8U)5<_C=f)f8H.aH
_[&)^,[GPK7PO\MO.d8\@6>UC4]cGI8cfe/E^>[K4?E[=&0K_G:OY\39#=Vd2I[3
TRWQYL8TWCPWGLGPf1^eSVYK32-=#GVcM&(bLD-Ue#-.N[0#/e-&6-0J2PgY)]H[
&JR/=]K?Wg/TX)QNb-#B.C@1W:P:P7TXF+Jg1=W8FH(\EL;.3U@](TUcZZXN/OXU
DF]L;F7FS1Q@[,aTM7eZH05O6#J7JX1W#R(?W(5@R7^/6_P/H=B0-PM4I;FgSC7U
0#LAf[a#5T1OLL2M4[O=YW6_M(KaS-61YY9(39\bEQ2_e,ZY20ENL.7M[&/XL+T)
gPXI85I(8LC(]UO&)+#aEg-@@10/I?T#)5^d6eO-PIC^)P4[6#DD/0g#,-[-c_S#
1EUEgJfL0:;B-Ub0f;3LB<J.,2#8J4(f@>.8V@I<H+f1)K3L>8@@Y6IXUM@,Lc(J
5S&:7FMbRJ?)YYbFS2H\_>H/P(P>b6^I-G(@1fJ(DF4?I/9#\Y[QI1.a2/A.BKQU
Q+ZQ^A)1(1T)3d;UTML3_aFgCJ6R\&E&AWRU.G)\))Zf@LG30g?U;a0(]=[OF9fX
,O22ZKRL;]I&ge)Z]/.W-OgPAO7=13P9\TQ-M>0X)J;&I&.G\g4g(0f0388LaI48
J2O7:BZY8V0;)=8EaUN5#LXLMYB4>R=K3@6A-UW;VVP=[(+9S+a3QbXgQ8M+a\I3
F42XFVA,a)Q9]>J4@+38=Xg_U;I4S;R\)_CI>&TgLB;;9dgXgH^K6eQ85B--[P-S
_I(>3+,5@bLBP&K2B(1YXNJ?.A[7FDD;K]P6QVKcO\>BI&:UG-U<8TdJdFgg<&-R
PN[40+FZ#QNX3D-@L/Te(>>^+,egP+-?W[U_/.CPF6<UVPL#YJc0Yd9eQG:\_RD)
K3KMPe9V\RdK[0D0-6V(JHd/#d0(_XQf/=0W2?dA>]4:]2)[=_@MR&9(Z@^?A1/\
M9X0Wc3F7NG7cffNRMEJIa&]LWBDO_@]dPIg7gfgO/ba-b#;.FY.6[^NR0OIHc;X
>SKL8[1<O_6>])FWBcJQ=&Kg,YUA152f5EVG6I\Zd4F\E6W?P=5>9ZGLX:3La):Q
5+Q.cD4T6T2gc<dc1/A73[2W9ZbZa+;=VcAG2X&>X3^dC:,5[C1O+7N-b^FfD(2-
^N]c).Z[aUa-SV?/QHOd[\1+Rf25;TTL:,7F7B>55/ZXHfBKdA_<QDgMC_@#X=Bd
UdE(H:BNc5c,[#d]-+RZa:P<GAL)3Y;:?)Bc(fZ=XaM[HLV@>@V0d2?Ug/)D-MI4
27:Y:gK<QBU=>K#U57,H>B+BB#Z>&7J,W5(\@?]JJ36;_QVYYG6GTG]+F/XQ_XgQ
FERCb@\@C9f26A^DCH[^FI-5Iee_)WBATTNF<gLVKKPeQ(034RH>^LVd4/aF:#-K
43&.7]_dQ&@D3-e^cE,1A4IKgD+6)#GURa&?Ne4YL8+&Td&d:K;_5=Jc3ZD&A.96
(B6<)7K.b-LK3&JMaNSAL+eD@WC]-EUSN);ERPeT^=8O<a[.A28V02FaY[JPAL4c
#>_A>g(f,:)BD4+KJTK921NHC3DDG,=Y\RX8Y<SG]@YJDZ;KD)F;W/^AZ2\BQ@Ed
)YX1[4<XM<]&;SZa4Z/J0:^=fb\dA?<5?+&02#N]:JG4K(;D7\H-<V4<=5#A+Y_Y
7Nb4NaaKT]I[1FR@[O\WZPgfA>&cOHI=0(A(2^Ae.X;3KgBK5cMRaS5GFZ,8+I)b
\_TV8A.JT/0Kf?Z>H_QbefdFcSa<]=N?H_:MRg[1JL)&QJC]:#HNFC#[\MA]8a@f
d>(Z4H#=&GTM)A))6,c3]^b\a^H&<W75VdCDY36252S>U;Z<>NO=\de#0E&K3I5c
I+d<\[0=33)A(0JgES<:PSK^DgCGKYd,+4^fHS_X;V-;g--K6XeDeKdRC=LIN9AA
M6]&UKM[HHNQ6/9])^JL:Hb3PZ<A3gD)fAERL6L_=b[bX-KYRa^d_d=-PBVQF>/g
SQe):eB(gH_@9b,SgJ-4<.+/MB;&a]ab+XXLg7T=\cd66(XAH/GN._8NcN/C?IL[
/2g@@8@O<YJ]3H_17V,?RK;0&-W0,=JRICgFZ(cEUNacU?E;R1JFA>W8+dX;GEK,
WL6Q]BD/22e_M-P0]KUM.NKZC4D/B(U,FQg.<B#G.<:SZ7KR#D>)050(</K@0IHW
3YaZ4[D[9+6<7<)c@38V.^1Qa8e8aHeZT1^3M/8:Jf[C]X9,fDea[N6abFZOPQcQ
9DTece6RA_d@Hg/<XP4gg,6c[Z<FT1XeMQ>52d1f]FKJ7O:3#Oe-63,YAR&[ZNR0
)-c(3.&D(YJ/[Z9O)Bc7#ZOa@Y:WB_KbXU-+8UbPb?CI+2GDS/E3<;bff@4H@E_=
K(L>_L:[&eV]-1H6=b)56]<4>W&=IIFMGdb1>8J1a),\<gF0\b3E;\Zeb-XGJ5&?
]2?4KUHd2^9QE;1PG&_1L1(=:3+P\R)]Zd.+eZHB8@G1.KgCQZ_U)EZTPG8\WZ>W
B]7M<;3CgZcQO;c>/FI#7AXadb-Z:ZYVbY8]NDOfUX^RYH7/Z:8B8SEE-c&O)4dd
M@d9@.e(\&I7@<K7KYJV,-DA8,PEZ3^M-)F7QcFJDXN,I=>KS[a1IaQ0:Q\b:-2B
+3YZ:^Ub.=[.Gf3QE_RHS:B=L9#JZB]JfcT.;LCK;)(aVYEGAb-I@XfEa1H.IRV=
[PeWOfB#X/dY&-dbFI()Q4T2e.F1DbWR9SWWM?)Y0PUT\K&(__6gA(Q./df?=cUc
J]c-C)Z515.=Qe>BWY>0W]g=+dGfDF&8O+e8:#4_CRVeA)I.@/]X);)=VU/gf26+
;P]&dKJO(@7B1:.^R/]>P0F2^(EKR_NTcFV\@GGFb+MV\MQBX.C@D+Ce9ZYN[9\?
=XR>=M2QYBXg;8M2KT[aD4I,5QS57[=UN+4GT7<,:b//=dM\FYJUA3+D(g70:V<T
OQ+KDJ<c2PGc]Jf/cV.gA6]O2AO;2#^FJ6UQXWgYJMM1N.fLY&V[IO-[E1\23:.+
BcJEOC_:IQ:E-^:f]7-V_b3C2b>d[FJLGUTQ&W--<_<1KELS^?A14[L8fS&@S0MI
O01:05#S=B)fDP;.Ec@eEQO=<FQMWHg^7>MZ8/2YG9MJKb^=0:c\bUf0AP@0?AGM
C9T[N0>HP_8K_[#74,YZ?7C?^:aI7a#G4Q[)-PD+<A4S&_E1:e4PZ.N:C3U)NC#T
+;bfC#M6BR2/?KAC/G6++[VJWFHg&-TU]Ub3+30I0XH=C4ZB#Wg6FeM+=EL:^PEL
BZU?>)S_OKgK##83?36T-Ee^/5O?7/9GOL[JVX:Z\2]NLMMSQ[ZbU@J9Ccf>JRXF
@9AIJ]&JK4/8[3_3[aCK1[QdE9c==J9UOa;OV^U)&H_F3Da9648W]IWT124N).UZ
::CGf\K6#&8ZfW-5GG8QKT,.HQ)fM;/^/:JZ;G@FN<.D?d7H;<JCBRfZ\#TE#Q-G
.b?=G8WYYab/]G5,@\fACXdIQ6(51X1GXBE?CTgdG>?90f2U),RT610gFQ<R?<]F
65^O1BOBaLLV/^II?@cGebaK.>?:4DS1Nd?M5UAGYIV0TD#UAH81SfTJ.D91RX,)
++U:\1@EHcg(?4F+I5fH:ZO62f(G6cX4R5[9I<WIf)4LC0PMSG[_82+2BIAKXI9[
cQKR,X]FN(/V)\X3KQc3CCU0Ya+6)[UTSE:Q(YAad6#.Y;Z+LfaQKC5K8=Cd5gK(
cJ6B<O)e\T2a6fgT/E/O7E6La_ATH/^EV,89LJQAWca\?=S5&J::R[>9<R)(@c[N
>7T,2BY53[;^eUc;W<XU?F+b>G6a0Q/L&>T&WGKQ<PI_@+M\.+^SB9F<]+XNc#:I
GUcU#LXe64\))GM\ZB5JV[B+@cFJOED_0^0_8[1G?62P0WCQ]>G9Da9V4@g.F)>=
.F2HN.gJI6M_2(N9e,6M7Z7-##YLVf83^TR;H#S[cfIPEQB42>;I073G&Y18:+W#
feOB-e@]JDGf/#NF)E+c2(TFWd:EO)3d@##@;a9I?O6YPCZ0YT,:=Z#G>BUaL9/\
#ZdKO.QG1e0U7A(57FE#=DaW51_^4<>,_Dbb=:2c32bR-QT9<4W1A6[)T<9@OZ;D
3?cXW;-^(?O^7D3(d25eJa,>041V7gTYGWZcZQ/6e=([:b8+C(1bB6N;c,;2D-QL
TAQSBg(<YM2W69ff;LJ<P^I[NQ:RYGd&g/?\PIQ6SFAXXZgX/DKW(R_]H,ETVN&f
.:>fc(3)IfQ]<H@[HH.E8X)0BU\R,8PQI4.WZIJcOe=W<a?+Fg;QON^N&SXgab@@
2\\JC:D8fB4fQR6@URA-)1IR?\)(7VW]:#]<I&\DHTT>eT;7b(Q0R,c,MI_51Fa)
9KX<RD]Q4bbNfe)TWbJ8@VdI_MOKDS[+F:\C[,2Se2V=HN5b(;cOMf&M-,?XYNPW
5W6RGGKL;L>S4WZa7aNKIU24)-8KI^ALZ+Hcg;RF;]QT@_71HL0,H45AS?,HG&L7
5I+1cJF4]<VaC60H&=;C&aD0REJ3MJK_A]b:/c=E+a#f5bUZcCDE4UbF\X]^YV&7
FYL3Df8QFN_/5>L,B;NdKC)B&GJ,&3#.O7S7.LTS^?314_1]E,4Nd0UUCJd\Q>\:
9;>fc+fIW];e3<[.X6J#Zd=/6ge=[ECgPe:^JUB0(;(RUYZ^12TbVaP7;QNBE6VL
1F2I:OL:=9[X62O<&bJMC<8:0;S^BE@ON=5OZ0?g9;GbT&5>H10X[[[.ZIZ^Q--g
[eXV.K7]U_C8K4g@[4g&ZV4_,Z6R(N\d0eWB#,dO6_;9G2?R8ZP?FQWI(N+,&KV5
FJTP:OVL((QEM=9SeYQf6&bR76&d<#.e:F83@e<-</gcG-+7@Kc:]6E(5+OT>9dP
dUQC?Z4MZIQ0]RT(D-PYbJ=5HHDTbg7744NfYaT5X42X7_4c/QA0^Y^c,MJ5W_G&
[K@MF4S.He7N#M\/#(V&R/gI5Ig#8A5bfd(<:.e(Z])>ZH3KM[5D4MGKa<SD?8Qd
/_?B+2]D4J6d\0&Y<YYIQSQ6_5-[7@[YbUE\XIOGJFD0JARG+S(.NMJ6D/L08H0)
E.6:_7Gc1LaHO]d913QZUYY#0/EU4UT^MN]C/cZVOc8>4eXKdbB)N^[;S]MMeOOU
\L?0MQYD4#;.fT:GPd8S8=-=UfT;IMQ?4F6VOVKMQ<OQXQ/]U/9G?/?6]V0#SBMX
3SJ4g1PE7X[dHIDNF@:C)3&C6&9,OGYe;1ZMcFVN&T/P:(eBb;VR-_e2DA;NV&/<
LS-X^HD45O^\,;H,DCd+c2^^08M:-Z;T^I3eN26>CQ?AX]YFNd@^?e(1FD0/Q)=(
V?&C?./b_C)-#3-E#I@927:3QNgAT2DT;EYa]<=EQP@E7#?;,?99J)(0eY7I,O_Q
^.@](BKd(7)P9g#IQg72^M9<@.KJ:P3C97JBLQ9KRObR/FLUdaE5J)XG\MWSV&_Z
::O&.Lad5a7_bT-)57T@4&05(IbW4H.+KOTCKTZ@\&)FG/Na3.;b7[QcgR(=/.CT
[>4c66^7IVcXPLJc?5Uc+MOJa4,XggNLQ54b\:A46gg#@7M:+6^b<_P_R^.bB..:
HAWKLR;N7VH6dSLfK4N+)dO]cec]YdW\IWQAT:R1=(-G1]4BAYWJ&KX>(:^F?FZF
,DMK-8ZF05KA8dAN;,H2fP4VF4Xe:>KADN>+ED.DZd1#[;-ZgC_[UI3_JC+T?W#E
#&+\cM4XAJV[,^@IOX(#32gDK4f#^5>LId<J#=-B+Ze9NCY1]JIb4aQ1(IZ](..]
30PN0.<TX=E+)2YRRJ(I:X[46a62;(]3b38&GWf5;)Yf#g_:e9c2V;TNa>:_\(<M
EZPg(6(7-c3fMOc?aXCZ4H]3<LeZ^dC8)Je3Nf=0(BQ+38FfD(c=Z2;Y99+KRJWO
f\07L+DW?+J<bCCXVa<NYG(dM.3+<;QSD@+Dd3KM05[=80<>(/cYFg,H.5;EYERE
0VXBSQ=[1CeMO>PJc+P_Y/B,G\?>7PR?44ef0LEg>,A.39ZQ\I>Y[G\BHRETNY:H
@TVe#N]RcK\4bNf=c:=.b769)YI(OM_-IeIJ7\TX6eSO0:Z(9?DC:=OcQGW-N-D.
H@P5Yg-QN#<CXRaG_<^CYdH@B^^CMI<gLB)CdFAU.;G=NR:=,N)G=eROWHH-J552
-231#YA,Y[&b2#\QE02bEPYXNK1?D(6W9SSZ]()FR^URY9W3[:>;8(8NV^>FFbP#
IP32&J<Wf.0#?6NEe);.#-X)L=-g,2#+]:eAY\\IYB>bM&d<&4^)VcaeN@eeID6/
IfY3N-.JDI>C=<S<)XUJF_XG13R92cdRBFeP?-D?Wd0aG.Kf9FL;.IW4?(],ROF-
5eN4WOP>;-N9_bN];<JS:VI=W,@V5^I0@YFG))VW7I12dfWO8SC#7W[C;HS0,LR<
[A_CR@U-4gPYB&^gR1=MX[^,\S@8)Y(^:#T0AHF.O(cSfE^(Ng_U#V(Z+?A0B6<b
J5Y<&#5<XZKIEY@NV&5YA-STNLGJ7AHK3S-cL0ZFe<VAS<7)CDK.^^V=6\(4f]2W
bKU]]PPRR7aRBAM:XKe8F/c0H]<NG@FU19J+9?_PKRg7_HVXXUNA-NI_VZ0_E(Ca
CQLN@eb()Y,PPD=IVSAW;Ncf9)?[FbK@9BYTab-bfO#&XHaG\a#HMP,<RJE1&4Mf
;MBJg.G;(1=KPOLFV?[50.bU<_R\Z_&RB9CG2G])L8(NWbNP&NGeW9WVd5e1#+=+
=,KP=Z9bG,S^.S&;A8A(1EF_:]deHf<9LC]+J(^J:Pa?SLFL@//PPCEB@4,B1N3Q
HJ9V>=2Z3(Xb<OZ.F[Z.IF,=;29_/EM(,&YB3>?CGE<,4aH)f<e#1^BXF&aeSc5O
(1g_;ZJ;?W@^\(JU>D2WM1ZZBSDA\WP6^/4RSHKGX+?E\_DXIId&-ZN.f,9)Oa+N
BYKQLH[@M_g#9O)_/bKT=c2Og[XFUe[QeA3@^N+Kf^I+#.JQ0^TEM22.de5U?adF
<8B?QG[,W]689WbZL:NFfW&O(WX_0BQ/U6K6.@,7DAU_5/TDaMT^.N,JPA7]^79C
B1[EHdE>G-2:2V=]1PV/U^F)YH;B,P=8_0]Y<>FNb?<,1/X3NFQ>NY<UKB>Nf+;M
<T/I#[3-NHe\,e>2LSXY6=R>cg.=ILOG546>NY^MZPNc6:>-5)L[[C=4KEbXPX;G
0EBM\G,VIe>;^12fJZ<M&DaMUK05>)fQ6F-X>FIPdG[.FS[VMDCO\LMC]W;/ZXI1
U)9O\&VP:6?B\ELY;e9egI<.=NA+7:+fdJ&Ea#,(Vf&2-C<#&dZP+7.O_31X)Q1:
?[1@e4,4K4:2O:6NUZf;ZH=DHB[\:CfY>YfK6I<GH[?B(/VK#F9A7Q?1a+]L(U<7
b__(FJ5DCBA5:](4c^N#-Z>9YbCK(S:J,f7ZZUJ;\eg6;T;YHC/Hb7FbP,48HJYc
.d>^/+O1(0H_FT(;Y-Q]Z:gPO,b_K@Q86>3B_^UDKb[F+,-&4#Ff8Q]=&1OH+CV=
_7W?9SPg[KR00E@gPKSCA8E50+9_]\\4ZcgDB:OP<e,THR24HUQ9F6Q6T\P#W1CH
>Ndg]<cBRUbI7G<2Z_.U+UZQKMHTUMMFEL5ZB8UF>BZ.gMgR)a>MHcR_:0->1)9X
ZZUS<I/Cb:c,-N.9K@UbV7[#X-3>]US<6d-I&O3ELfOUe^S-EVR+[H,F]3FDDMUZ
f2:O=H&e#I^2]T;80?g?#>dXT&<B5BNGG>)9@^2\O2:0?^T6b]+^(?)>YS_X[VIa
cS+(dB+3@]NWS5a<QbTf8AJB,WW.F@\1=G3E?_:>AA?>,Ha\Q0<MYc2[U4:75-UH
;@@5SP#:Z-gbd>9(EL(b\E7U.,K?7B5R2)Y+?)5L>4:bA4;M,PKTX)+Ag)<)J_4C
a&I<BJ);<38^2SYZF]HG11D6\eU>g8(<CfH<^K[Tg^SM5OH:I3SfIV7gB:5,ac3Z
QV>X+/f(10>C:8bHc-CZPZNFLfXEE;ID,H-cJBGgXb9NYBFUSKJW-5JOF&Yd)g\a
\Mg8g(@_NV).95UMRL7AeRJ7L0\SS(Cf-ZN1=Y;7)#cd;YMWG,7<=YE)H)+MJ4,K
Z&>7.\5G#-LBG#<&D:F4egTc^SNa>_F7-)01V+VF=2ZX/FBgNN&,J_:>WDEYXC;3
a:>+JTC6?G/36eE-_[cF=?E\.9ROGWMYf8ND)QUMJT+GYfc@DWJHLeICK9<>,\&/
]6:0#LGF)\]M?;6CA:^YH9N?:9-eHL;X[IS<eM//f^ZDSD@fe^W_U;GLD\\S8PJf
B:6B+[W/ZM]=<KMPE;RR(C]6ZB.?\g\TZdJQ_&a\Y)#[Z=&Z(0Ff[HEY05egaJ/R
56Rb]0X/ebTH\>H_aGYEU-:Wa.SI^BN5@.S?_DN:a4a[Rb3.N15\^TX,g?L<0X(8
9[[2(TS=AW+5>d=+[ZdU^V:d,+bFTIcK5P>BEa4Cb#D0R9V0X##cgSMA_/V[X9WE
a.TBIgLX]/R#=g\-(+EbK9Z,OSaG-PcF?B27R-J:Zf^2)cO=ZKC4=>4AG-0M6AJ9
TK3I#2)_Jc@efa1F4O<gc0\(\&5Na3#)XG7/T163]3<D36,DFZL,Aa/]^d_-1]\R
XM[_+2L/>?,SdHQ\Y?f879P3^-/RV#6K=98T49+Y.1JJPU08Kb<7KfGF&bR49LD3
RAJGgWT/,;Y+IgJ_)YD7;>[S?12^6>L04;60TgKP?gEBQI6BDCPL&6#-JEcf.WOP
0UdPXU40AET[]0#4?&M]?,YS+13\9R\8If#Mg+-(TD9>=_BX\eTRf4KeBb65^>O;
\PV6CbfH[IR?cVS_F?F&Y&E_DGP+CHXVR>[[[Y_9XRE;,#<JB;:(.N7>EB^FC/]H
_4dI4O_+F65U-L,KV\F(T.,+QP&)de/W\?=Y(KH/ZRa(;\EB@6+]CReZD&.N^a[B
M?dL_3&eBR70)-P_<bGc@5^SHUS^C>bYN7eTM/KG1+T5W>79G9S&L;XOaE3.B60X
_OPMD/MSF832Y#R-Cg0.H,/AEgd=B(_/HILX[<?d:eP)_S7)-dJWG#7,N6_I)GF.
g1GgLe^2YUJ53Z#40VcNET17=TYOA]a@#;TH5VIFV\f2E..<5,G?]5?Wa5Zc4dCW
ESZ>7:=Cd,,P[6e1#4MN-VQ45T<.Y+/)LdL=PTa,/-49RXQJ6<?^]-4,WE?Sec)H
OW]LF_<:3=54GR&HUY1OKLW@W@&U5/_?97QXe]V)_Jg1530BX:BI[O;)AAE1EAeD
1gAGcRPMJBd7MCeX>RU/.GK4A3963,1^_CJGZNL[[H4;BMLeZcb7[G(3Sg?/AQCa
aK^M]7<:0=R/J:c+:4X[/WFBN3DLL(:_SXW[L^MLGD:OQ]0a3Y)JIg9ISWdd;c0P
R;W8.J&KGfeDaR=(_bISH7[PA:cXB</.Q@(ABX\5f<U0:7(gS:.V1:e/NM>V]17A
3ZE18;f>Wf,R1?5:+d1YGTDMNKFZC-fR.\C7,LGAM79+057A]1d=GdG3e/+7;FMU
If(LbVMYJ8c@6ZXCQ>S6dF<T>KM-LC-DF?:9)eDbgUC>N3M.aI\feH1g2bCgJPTd
-P:;b8HE7+cC-H)7CN-.[:=U)@5@:Jb:D1?9HBLIb&LR=U_9[>I>M:C.3#a2<UZ]
D[]<2d/]\WAC4Z8GU-@<Ra?,U;U+dDS7O<(<Y[O?I#T,TV#^cXU=G09<U-W:K1f)
3S0Hc+]TSJ0?1HA7e#DAY9W@4WE_aO)eJ]R870;9&ZIC\?IQPTA<HV?D_#QeD&:F
HY+H+00Y0]U=Gb]OZ3EDGW;SE-8X-])_V7Y\2&.=[W8YdZN@1g\dS)Y\+I];IE)7
-7eA)931T&a8NKS0aPOJ&7C:cY,Y<+R.<RF3;BUQ/4\8RY@+;#2Gd)5-FY&TD4^P
].M[G+4^6Ma[S^G\(,?:IPQS;N[9YPS7AJe3D&-<92e0B=fM5FJ?5VMEH+].41/d
VNV;#R5@eg(OCfIMF\BZ(SUe7d)4C@-1O.?.fD?IdR>_1Q_fT1#A8g90b-;ZY@4^
DPND?_E9TM<>3K8-44U1-@)1;0T/5LgdZX@#+L6H7)4<-N:XeHJI7<ID@cH6:&_Z
g8&M&\bCK;Ob4K3R=ZZKW:2_<,[PV@Mc0,P6J\8U3H/<YcM2K8#.JbPMDT,XI\E<
J<98UY-VdMGE:G;7K7/O14<e<X]Y/(28=Q&?:YFUW;C+,:SEc8#g.XG?M>S8aUA)
;EJB7Ga=IK)Y:OO(dUaPJT40SDE@\P(;=fba_Y\#6KY/CFR3JGH?G/J@J2_-bU)6
+JfU/=[,P,#)=>./X#5]I7+=c++7/#D^(?OQ+A1>P65RIDN6W,^Y\>OCEa?5UYe4
5V6b4[TQD2dKRdDN8.#/9OKS)_[AcdO[KVF:5aEd\O#I95#Se1CdSL?0c=M.(FL^
YOR6+gLAMc^_KMTN#DR9;Z>ERf9:=O1V)4_J5;#P&HA&#XPL0A=55L[\@Z4W?AJZ
f>CWe):dP?ZQ[4[Q-QAEPDCeNBdS9F&/IY=7F@7,25<V&c6&-Ra^0cc90P63?D,X
e4.ULZ.A@DS1eA^N6]@BFHXIMaM@6#ME5d;NEEL3[JUOI1Q7@L:)4.2HD)UgFDE@
KXQJSUQ7c9\2O^bJ4=&SH8&If-#E;Q])9\A=]VB.+P_49_+f^BC)ZAGLRPW8\d/O
,8VGFWV+::A#e1>T==2<IO1E]@8Z&0SP.eS8)&)YJ,B)S2.:aWE77/XE-<f1:R2#
\2RPNb0DX>0O=N>-YTOV9J_<39=LgT<B_WeRJ-^<K8\])H>S+b53g_S+Od@51VS/
dABB:bNF4/+068f-5:L6dLAZ(E2-/LQ,W3>L9DW:8+^VD2O]Q_B2-T6>MCR;_7JX
/eOX)=S>Q7C>@>)N)IaJdeN#RM1?_g2[7bTRTe7<V_g)[>9K7\)H@Lbd9D5cbSJ3
T&JQPBG(:,\<W;;eV:;U/2@8aXBJ;^[+/#KL#0+E#C.]I\9#Tdc6@0X?<<g1Q8W9
QTP]G6>)gKG<;FV-g+bQbDTc_RED-C<1>ENA^WD1a@\](SGa>S\/6OZMWP/B5K,W
8D.1:A3U\&L--BA7BJ>)KKD7A6LK9O[O[9N=V-O)^(X9>7=S=/>L@1[;gg_3CE-5
RcM^VY;:>L=HI[C3d12I?ELN^U):L<0dKegYLVcV5VM_6Z[c=+/JKFWS;?2O#?Z-
GdN:La+F:YGe95LSR.NeJ9@/R4T;Q9I#JdM2b[QV#8Y]YW;<WJAN^8;..,)<Z89W
PRA.@g\4C6NE]FP-T)@009@<LYd#bT&70ebVMQ++bdc(5C3Q.?GFJ+D)(5UZNW-T
@94JJaf.DKA\T,4HZXLcX7=2==&]N^BgeOT3KKZIc+K<E@BL6,_FdG8d2K(&g_LQ
\EVTARd<NK/JB:RM5#TN:fP6+,XE/d;6F(BGe0//IX5)W>&gY^9J5+W03[Y;d&dW
U-;/7A4QVM@_]PHAS>cW9b?<edeLS^bY6@)C<O&8T)F/U=U>S+8XXFe^?\T]]a?>
TJFC9AbV[c8,C.9JfM0:EI(-Ig)GFR[Q)IRX5&b7ZZ[?VST.P=X>TeV-)&;/aWY^
UX]_>@:K39Z3]&1Y8ADVJX;VK71Z+R&;1>\H]OHgfgWB-XYOYc9VQ#EK_WC(CM13
ZV72KgQ/gGdcA;,gbR#gK84#Vf3d4]2;GBM)B3bNVJJ66Q+C>0GMMD8_8SCWe[Mg
ge1/1g56W7GbA:;<WC7LMed8<.C-YN0SC_cD)@<;+\\9^.],;Z79:+FQK0QVS?>B
&IY82a<W5;YQ_#bRR7(UcL\Q+J?&I_R5,752U(0).4L4C1L//MW.3]Z8f3A.Ic7B
HfZTCPTIBXKU<4,:,NTFNfC#B93f^I?_2A2/(US6=+2>G5D/&R2\AD.NP/N]YXg:
8RcIgT,:F2.:UE&S]K<CB3GgB-6BDcE<Q?3a74b6VaaPc_/Y9C?E\1\d,;^dbdX=
?fADBJc(FWAa,5B6b3/1AE)&R_#a0IVR9e]YaLdKVDaZEN?aYa9284R&?YgZWV6)
)=E3]NX\[L;5B^:SU&?)fa)&7:WdD[+MS;;OZIVG#(,cMg>-6ZG9#>Y<ESe,RIg;
#T4f7++HCYPgRATCX8:7(/55_TUg/Z/70R7g]#79T95O+J.3Y?a7McXYL/?0[4dY
Af0c4/2gED/ZZY@#9&B7HKA0Gc@Kc?LRZ^^VVb8R?47d0VUYb+70A;>)GbO#L0MB
8M9gQ_>MU[BT^UcO\GB[(FZcVE-2:#R,23>[H?FA-2CP>VIKU@I&1_9_6YINb2SA
AI+9=CZ&aQGJDE;^(C6Eb(+MPXPM1VfVSb1[7A?aC2LVA[V[JUV04<BPF3>H;LU.
b6fIK7(&T@d3Y7Y,MacLAJ[)&-f+Wg/:L0&-/A@WaIPa^B80K9Z0gXK=@?IVg/Ef
Ea=TV\6RGSM(N_O5&f]d\D_HRNY-fPd-Y?Bc;JHa<#T3^7AWHfQ@W77E&Q6?I5]?
F<-JL9-Q;XS,G().K;/S0AWC.K4ab\U:L=RO7B&3O32(X\]<f829-HUM+/1+CZ.U
e8aZ8/<9LB/_#W;_f>7f2Ve>PK6a7f?[\WbTUdX7Df4_faSPaHF38;HU]ea7e;/d
M;LEWS77PT#]^<.=^EYU25L/AH?&F;9[J]_BV;KG@;\Z<[OWPOfNA59T&?)7QWeS
2CG\>YZJ6_1be)VR5cH;G&<eL)^gfVO@?dOd)ZW)2>1\BU,J#,/75H8]^#?))LIB
2HD.d:S.;BX9=#JD/PIcI,^.1PFF\/eGfTT^V]]FG=JDGeJ]<TU3CA?QKLF[YPd^
S_-a0b]0eP1^G8g>KVe-bO[CcXBA@XPe6ZJ2RZS=7.Lf\N]QERBGO0,NZ,&[J#M2
aY_?+S)O+1&QIF;)F?WA3Y)CP0EB0WD:H:<Y+VRS157)ZX>MV4))U--d0FY+K;N]
(_M/D-&W_G7_>H2IeKZYBBSUCE()-4G/ZZX5,_GgaaKO:^<^/=),-_,:(J(U\8?_
7R^)?(3UQcTKR2b^CcFC86B<I1DA+6(4Z-G1Ea6]POP^c0FLJS9Yf^F2/PINLYW+
]-8T9?J:T,V_?.Y2C?6+E7;[:=:K^(M#>ZK_IW7(/]>1R;8\VZETY0Z8JJ:AcH9d
MfEE:SXBeQf^cJ,/2W:ac&)90(-\#A^b[EcYJQ.C+cR;::.QT65@d-5;>Q7]]5eJ
&HYfVE(.>-U:b-W,KWc&A4L]b>0W?6T-[RPXG@K=2.BU&,T+ea7If2/N2J;3a-5>
8/M5CCW>ZRZ+c=A_3]N)4^ZXS=b=--.bR+]<>E0=6B8EO.1BJ=V9+3V-V<G)#Q8\
dHFTT_JX7Q[U34KeKX\Q^HL1<XPgcV,dO^+]5\9:OAc?fKR/-H2,/@J.c5JV?G^?
,HXQ4J)=6>ce&8)SGF]/EcC@XD;FZ]CaD6S?bV5ZXB+6Ue8E]-Y/f2MB7O8;.<fC
P&U][e^Qb4)K(8@IPgM>-b3.JF-J]4KV3TP(EVY?K]IEfaQgWBKLU.VR..<d7eXa
[=.^<,<C8X)\<EC:G44QL_OLV)e:P)65M0]8Qf60gIV[IX\<M-YFAg=3]#Na@(Ma
N@EY8Tf=>PTCG.-]B91>bXHZ&X0cQYRC2BeI?c-]aHff)#3He.aA1PYf0269>#b5
O+P7V0@\1.YKB/[W_&_bE8YLL08OLIP1Y:IC)X<^4M)1:>BY5A([gG7:E[SXS_@[
OA+VP<K(K(;a5d87P-H]W03]@7Cef1bW3I)(G3b,7(\Yb(_JWQD>5^gLSM1E4C8R
THGa2RJ9Ma]S8T6ccbOEQXXgcZ;8a>Ed7N99\eSB[&bW-g<(bbUM#_L1aML==\dM
6#0VL9&4KP&E1F@A+Z9c=(<B.LY37L)BG1M<Q-EU4eG-K;fNX[8.,6E0dWV0Nf4P
2>6-LP3;Xe5RI(7_MZ[>&HZ>d#@CG\.(-QLK>MgMOCN4@;^cdAV+:<MJM5MR>,([
[R6TV@&>3J\>ETdeAXeT:gN/AT#UMAN7>B0W(fSY@e47HZ]H4aJ,LMC=D2M)<_:J
L8EW4@&:V(^3#/2b5GZ6dC.=.?)L#C(HdNWZb8&I+](eS^?AS8&b#C34dTZE8M29
D,b19T<]QE@7ODT=<EI+L/^f;L(IeW61c3K3H57.\bJc2c.NH+Y-fcA],PB7=aU8
_+C-U7B@;/_)^=#^5#RA1G?aO8A;Q&/1Q_QbZ>.7C^[1I0@b?-L@UB?[GHH7aCF)
TJ?>Y(dV^^GB?Da(HL\S(ID@?E9W<1#S2V7<-)f[XS1eM=(E>\A97T?^N9VDOXe7
D+<LfAgRB(0/N&5Ea-L=&R;OLSTVBZ44TfC@K?UAMQ2Xa0Ee/E(a]@6b9IJ8aSce
#C8g?bB?95;;\eHB.bb_#XS0A&a(O=#D9If3O4ZX6fQ471J7a=dbd9HP6e(2(.84
[U/FEMgS_A[+;bDBL<)<WI8UcV=;+g/<]_&Bg(V#D&b]bbXG007Ge_.\3XAg<GHW
Q,+QH4VB8>=U90S\PNd<25]C5EF:8:Z<L&8,R3K@Q,(B)140&UaX7N<_0)5.9DgM
O#-CIK26CGg,SDfG46A(aM1@X[Ye3;9LZ(56([@eFc;(6Cc90&a<0RYef2H>H<fg
-3Y?[^GaOG,#A):WdQ#3:,SP6QZ/@I6NSHLFI:G#G>&?;6[9X=W)&>_Y6b<EH+.>
ZX5PNT=#;(-.K2O.Q+J.^5(^5RTZb?ZaIM;GGeYF-TBWPR;GDM-;])0Q1USP?9&<
ALc@W1=OW<??d_#)4],3M^SKXQ?B5[X:]R>R2(W\G.YR@?4T#c\J1bd(_(L3KWN>
JfeE-dd-UH&c75JGE)SVAV?A?-Ga,\5MQ?7DG)+([(>#W7_9MT(>HZ2L2)a/5\5=
K0-e5S/>b2\FKCEHNI2B;J>;3AZ&5,Mf)#,-=VS<KNI=&QH\D?++G31E_dTPd=>U
3&C:U6V_>60.2R-&G/6?8+M^.WVAYSH4E,@#_K)AOEd?b]_,A.PfbG]Db6Z0,(a\
RSQ,Bd34\EU:?Qb9\S74PPD1-:R/\](8,gWc+^&d1OW3?dA+Ofc<fcJ8(beVZ=BV
7OIA^MfUCY8PU<-Ig_51eT>_M++/&ZY-H/0.8eCe^&GL+A+5H?83ffQ[IKEf14Y&
eLCfWcWOF0]G0EF;R(>]<gIbCFcH,O(9ID2^+3FaCd\)B4.&+Lc<f_??KgO-4LD.
H67JSE+JV_MF1-_50JbSe;NGQH<T468B_FJCJ7CK71(IWFZN8^P=:?S5)&H\VbfK
QN9TXGcU/<<U5#5eVX7?L3M/gX&gV(X\=c<&W9<b8e0OT.a<M2-dQgL@GeQ\a2-H
QCTe)8_OKE&fP9LdEOWP?EQ3?Ba#3d307O[(5,f0R+[O/SYC5Rc^/V]32W0_2,+d
K-]F>F=UL)U2\4:Jg37Q:G\;IW\X_TNQ1BAVEVFT+86AFJ\E79CIO]0F;#C0WfX1
b1_DO?2_I4A80<S,?Y3U03/d@PVTS1d[(K=2_R+QTgEZO<#0\LWGJFO;=2V@JDe1
&=[6USU:RKQO6,^Yb-Fd5Pb:HLVNBabc,8[X0T3JU0f(S@\@&WAF)\1SfQNJ-;^5
G8+BIO5;@ZDOfaEG4M4@_8Y^_e(?Fe))&AJ6b@)9I#D2S\DcFbY6PecP7dBeEWgQ
+56,=>5ZI-Q38F<V1V/Y&N,/g+3O3:=<,8(1G=>HS.B0>^TCCf^RG:,^R5Lf47,D
48K1[5?3f=R?cF/>eM-()=JBC5.7OFK4Ab=I\VT0[F#C;#M&fdgQeL?.18UW0RP[
]6KBe89^>LI^PXG:>L16A56R^ff_F81:WcNF(5&JCZ=a3?=;E]]O22()>=>Cd])S
#bXg]gJO.//^Y)^:egd,]+1d81NNfa@e,#<_\e_5Z7EPSM0_V)P9897_e7VR@5-O
6fA_eM4/]2@;)R0b.8.N;Ff_YS?N@1-NW&c81.A9+LV8YJ4F@eOC4ASIM41Ab9=.
RY^JIeRR][/F3F(/Bca50@a64Q1)/-/<4Z[gdcd\2S]c?11GM;[>X6MbgO,f.P4K
F5]-XXK2L@+[?LY_(#N/RM;b(MO-;_7A&ZMHKEJ84BW))1[33EJ8DYfT7>,=(17+
M<#VbD;F6I/[@#b/E;UMJE0FBC+NY?>2W<&)2+U/8VGMXDQ0?bW:FHFD7A7dL8eL
6A](_G,U_GSMO8cC>S0gCTK-LJOaM+6]TASL<.80KA<]&E7aNOW2feCMC/RRJSX5
R(;7;60\cSSB)5EX47.VNWQY002Pb(GW&PU-ZQ^Wf0\9-:8HHec]T,76@2\=aC9<
6<7:B-W/+aR61e[X/C\JS-YEE1IG^@LLUFeC&BIXAY]<Ec[BSQgaM_<_</;PXYJ3
/,0LP8\\&7S&T/cA6SBG-3A,g?#/U43Mf0Y@)3QbeHBZ:6J#M?0\D<ZTBb)NP>f6
Q2N&O>cJAe,SX.7>X2WV6Ae;gFV=H;<b[:,O+EbC846(PS:>8<8OEW;9G8EOI\9N
b)Q)UAb#(<<[,Zf_@4@#=:=E.Y\;ZK1N(g6.59/Q[XU67_R]9bO8L8A/SL9JI5?C
Z#\BgX6Jf[e>]<(0\8IcWD29NVY<-0M@_H(#U]WZ85IMI+N@F:U+FM6a\&)=(.=\
NE5Y^386#<NgPQeOT_H<PQ=]J;==84];bYW[&3.fM@IG=A.+Lc_+0U_=M7C-+,+B
O48#beCbEcL#J2LU\eT].1c7eVV06R:>X1.[K1dU0@-+DV+(^U]g^Z2M]a\M_U;8
.4b((_W2[0HeNZK#>CW2CfeDQ7_7M8(I_^)NaEL#)GMf1KTJI^+T7U42PKJ(SU@V
95IC+C76VLaHF:G&>KM@#Q\fR=8OO:=-?E#3BZfL.gb/J6R9&^DQM/_T;R809E=#
Bd_#I22,3F&Q@SKd9AS.6+]:U:a44(47a.,J.Xg\2\e;#aG_cf8QFFe/gAGD-X8f
W@?QIA29RJ2P5NZ5cdCJdHA8-:-2U-WO6/?_/d(_P]W8H=Ya9SaA.V@VW_-X]6[#
?d#&\=E]#3>JIS+[2]]6MZI?(URG-c..cfAPV_GU7TL.-5=KZQbOKHE24OQ+bbL(
G#<@UM9P#d\]\Z#-NP.29Pg3WObTD-OJ1IJN/Dc^?0\a;;Zd95Q^J[KV/fF^FF;3
+Vf@_)bKYfML:3fA^&#+YM)dII^7.P<f-2H98MG0W(c6bMf/49\fE(T75=5Mgc1D
@\:8cM2c?7_=O&@W]9P):>9eJ<^M4_V4g4PVK4I/D1UADSBe2b2TcE7gGF-]TeWC
>>a0J62U3<5F)0:CY2T9,5Q[B;7?bI[@@^GSX[g0\e1gQCXK1<P:PCc:_2e.Sg;V
LRX0I7Lb;&bZ;eS2Q2]P1U6O]:OHfT6Y]<.ALQEPD-U<^3<K1<>@6L>Kc)JQ-NX+
S;IG+-_P8=gbb5/-><+DW\9/W5=),?3G[_&BU<0S<G[K:61Xc@H_Y7[8\DU875ab
GMEbg?J=8ES@H?cf,&8M?2VXcV)J0(+T[)4cMCd<+.HeG8KfeF49FBH-f34gWLPa
\UfYI(?WeQf&?HM3ZS\eEaGC6K-4-KP[ZR;84@F;3_Cc7IY-.14&[K:CK#9SQ4IY
;/LWGZN(EP0A-#YOLO,,7c6/7+#R[:(_(M;4UP1D<[f#F<YW(@eBL?f(-;+eQdbX
NM73\1>;J8SdVZOHVO8#d+-\IZ(0J1PQX66XZ_[]?,\XMXA+I#YAP\-CcFDHN3=^
90JRB>c]_/?._>^7IabdZO^5Se].:Y8EF(RNT6Q]Y4RfF>.>b3>#Pd_</9P&d#I(
@LFg]Z#5U>[=]MNTXa334;(RO#O?H)B6^3TC9_G&8K.K+Q-JM7eGYQ#b;9XJe;f9
.O1W-Ga5<WDJaYgR_.8X0RES2a^ESIaXgKA0>.=X589D1(f)5<OF9[IffdBV#,Q4
HOeX(K5.a0R_-Md+\>\(f<R=U(AG,Y\FdPMCOeE&f2a&R+-HReP=QR0AE21[O.Q7R$
`endprotected
endmodule